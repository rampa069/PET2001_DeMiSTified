library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"741ec04b",
     1 => x"87c702ab",
     2 => x"c048a6c4",
     3 => x"c487c578",
     4 => x"78c148a6",
     5 => x"731e66c4",
     6 => x"87dfee49",
     7 => x"e0c086c8",
     8 => x"87efef49",
     9 => x"6a4aa5c4",
    10 => x"87f0f049",
    11 => x"cb87c6f1",
    12 => x"c883c185",
    13 => x"ff04abb7",
    14 => x"262687c7",
    15 => x"264c264d",
    16 => x"1e4f264b",
    17 => x"f4c24a71",
    18 => x"f4c25acd",
    19 => x"78c748cd",
    20 => x"87ddfe49",
    21 => x"731e4f26",
    22 => x"c04a711e",
    23 => x"d303aab7",
    24 => x"d3cfc287",
    25 => x"87c405bf",
    26 => x"87c24bc1",
    27 => x"cfc24bc0",
    28 => x"87c45bd7",
    29 => x"5ad7cfc2",
    30 => x"bfd3cfc2",
    31 => x"c19ac14a",
    32 => x"ec49a2c0",
    33 => x"48fc87e8",
    34 => x"bfd3cfc2",
    35 => x"87effe78",
    36 => x"c44a711e",
    37 => x"49721e66",
    38 => x"2687f9ea",
    39 => x"711e4f26",
    40 => x"48d4ff4a",
    41 => x"ff78ffc3",
    42 => x"e1c048d0",
    43 => x"48d4ff78",
    44 => x"497278c1",
    45 => x"787131c4",
    46 => x"c048d0ff",
    47 => x"4f2678e0",
    48 => x"d3cfc21e",
    49 => x"cbda49bf",
    50 => x"c1f4c287",
    51 => x"78bfe848",
    52 => x"48fdf3c2",
    53 => x"c278bfec",
    54 => x"4abfc1f4",
    55 => x"99ffc349",
    56 => x"722ab7c8",
    57 => x"c2b07148",
    58 => x"2658c9f4",
    59 => x"5b5e0e4f",
    60 => x"710e5d5c",
    61 => x"87c8ff4b",
    62 => x"48fcf3c2",
    63 => x"497350c0",
    64 => x"7087eee6",
    65 => x"9cc24c49",
    66 => x"cb49eecb",
    67 => x"497087cd",
    68 => x"fcf3c24d",
    69 => x"c105bf97",
    70 => x"66d087e2",
    71 => x"c5f4c249",
    72 => x"d60599bf",
    73 => x"4966d487",
    74 => x"bffdf3c2",
    75 => x"87cb0599",
    76 => x"fce54973",
    77 => x"02987087",
    78 => x"c187c1c1",
    79 => x"87c0fe4c",
    80 => x"e2ca4975",
    81 => x"02987087",
    82 => x"f3c287c6",
    83 => x"50c148fc",
    84 => x"97fcf3c2",
    85 => x"e3c005bf",
    86 => x"c5f4c287",
    87 => x"66d049bf",
    88 => x"d6ff0599",
    89 => x"fdf3c287",
    90 => x"66d449bf",
    91 => x"caff0599",
    92 => x"e4497387",
    93 => x"987087fb",
    94 => x"87fffe05",
    95 => x"fafa4874",
    96 => x"5b5e0e87",
    97 => x"f80e5d5c",
    98 => x"4c4dc086",
    99 => x"c47ebfec",
   100 => x"f4c248a6",
   101 => x"c178bfc9",
   102 => x"c71ec01e",
   103 => x"87cdfd49",
   104 => x"987086c8",
   105 => x"ff87cd02",
   106 => x"87eafa49",
   107 => x"e349dac1",
   108 => x"4dc187ff",
   109 => x"97fcf3c2",
   110 => x"87cf02bf",
   111 => x"bfcbcfc2",
   112 => x"c2b9c149",
   113 => x"7159cfcf",
   114 => x"c287d3fb",
   115 => x"4bbfc1f4",
   116 => x"bfd3cfc2",
   117 => x"87e9c005",
   118 => x"e349fdc3",
   119 => x"fac387d3",
   120 => x"87cde349",
   121 => x"ffc34973",
   122 => x"c01e7199",
   123 => x"87e0fa49",
   124 => x"b7c84973",
   125 => x"c11e7129",
   126 => x"87d4fa49",
   127 => x"f4c586c8",
   128 => x"c5f4c287",
   129 => x"029b4bbf",
   130 => x"cfc287dd",
   131 => x"c749bfcf",
   132 => x"987087d5",
   133 => x"c087c405",
   134 => x"c287d24b",
   135 => x"fac649e0",
   136 => x"d3cfc287",
   137 => x"c287c658",
   138 => x"c048cfcf",
   139 => x"c2497378",
   140 => x"87cd0599",
   141 => x"e149ebc3",
   142 => x"497087f7",
   143 => x"c20299c2",
   144 => x"734cfb87",
   145 => x"0599c149",
   146 => x"f4c387cd",
   147 => x"87e1e149",
   148 => x"99c24970",
   149 => x"fa87c202",
   150 => x"c849734c",
   151 => x"87cd0599",
   152 => x"e149f5c3",
   153 => x"497087cb",
   154 => x"d50299c2",
   155 => x"cdf4c287",
   156 => x"87ca02bf",
   157 => x"c288c148",
   158 => x"c058d1f4",
   159 => x"4cff87c2",
   160 => x"49734dc1",
   161 => x"cd0599c4",
   162 => x"49f2c387",
   163 => x"7087e2e0",
   164 => x"0299c249",
   165 => x"f4c287dc",
   166 => x"487ebfcd",
   167 => x"03a8b7c7",
   168 => x"6e87cbc0",
   169 => x"c280c148",
   170 => x"c058d1f4",
   171 => x"4cfe87c2",
   172 => x"fdc34dc1",
   173 => x"f8dfff49",
   174 => x"c2497087",
   175 => x"87d50299",
   176 => x"bfcdf4c2",
   177 => x"87c9c002",
   178 => x"48cdf4c2",
   179 => x"c2c078c0",
   180 => x"c14cfd87",
   181 => x"49fac34d",
   182 => x"87d5dfff",
   183 => x"99c24970",
   184 => x"87d9c002",
   185 => x"bfcdf4c2",
   186 => x"a8b7c748",
   187 => x"87c9c003",
   188 => x"48cdf4c2",
   189 => x"c2c078c7",
   190 => x"c14cfc87",
   191 => x"acb7c04d",
   192 => x"87d3c003",
   193 => x"c14866c4",
   194 => x"7e7080d8",
   195 => x"c002bf6e",
   196 => x"744b87c5",
   197 => x"c00f7349",
   198 => x"1ef0c31e",
   199 => x"f749dac1",
   200 => x"86c887cb",
   201 => x"c0029870",
   202 => x"f4c287d8",
   203 => x"6e7ebfcd",
   204 => x"c491cb49",
   205 => x"82714a66",
   206 => x"c5c0026a",
   207 => x"496e4b87",
   208 => x"9d750f73",
   209 => x"87c8c002",
   210 => x"bfcdf4c2",
   211 => x"87e1f249",
   212 => x"bfd7cfc2",
   213 => x"87ddc002",
   214 => x"87cbc249",
   215 => x"c0029870",
   216 => x"f4c287d3",
   217 => x"f249bfcd",
   218 => x"49c087c7",
   219 => x"c287e7f3",
   220 => x"c048d7cf",
   221 => x"f38ef878",
   222 => x"5e0e87c1",
   223 => x"0e5d5c5b",
   224 => x"c24c711e",
   225 => x"49bfc9f4",
   226 => x"4da1cdc1",
   227 => x"6981d1c1",
   228 => x"029c747e",
   229 => x"a5c487cf",
   230 => x"c27b744b",
   231 => x"49bfc9f4",
   232 => x"6e87e0f2",
   233 => x"059c747b",
   234 => x"4bc087c4",
   235 => x"4bc187c2",
   236 => x"e1f24973",
   237 => x"0266d487",
   238 => x"de4987c7",
   239 => x"c24a7087",
   240 => x"c24ac087",
   241 => x"265adbcf",
   242 => x"0087f0f1",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"1e000000",
   247 => x"c8ff4a71",
   248 => x"a17249bf",
   249 => x"1e4f2648",
   250 => x"89bfc8ff",
   251 => x"c0c0c0fe",
   252 => x"01a9c0c0",
   253 => x"4ac087c4",
   254 => x"4ac187c2",
   255 => x"4f264872",
   256 => x"dcd3ff1e",
   257 => x"4966c487",
   258 => x"0299c0c2",
   259 => x"e0c387cd",
   260 => x"def3c21e",
   261 => x"ebd4ff49",
   262 => x"c486c487",
   263 => x"c0c44966",
   264 => x"87cd0299",
   265 => x"c21ef0c3",
   266 => x"ff49def3",
   267 => x"c487d5d4",
   268 => x"4966c486",
   269 => x"7199ffc1",
   270 => x"def3c21e",
   271 => x"c3d4ff49",
   272 => x"d4d2ff87",
   273 => x"4f262687",
   274 => x"5c5b5e0e",
   275 => x"dcff0e5d",
   276 => x"c27ec086",
   277 => x"49bfd5f4",
   278 => x"1e7181c2",
   279 => x"4ac61e72",
   280 => x"87c7f2fd",
   281 => x"4a264871",
   282 => x"a6c84926",
   283 => x"d5f4c258",
   284 => x"81c449bf",
   285 => x"1e721e71",
   286 => x"f1fd4ac6",
   287 => x"487187ed",
   288 => x"49264a26",
   289 => x"c258a6cc",
   290 => x"49bfeedc",
   291 => x"7087d8fd",
   292 => x"ceca0298",
   293 => x"49e0c087",
   294 => x"7087c0fd",
   295 => x"f2dcc249",
   296 => x"744cc059",
   297 => x"fe91c449",
   298 => x"4a6981d0",
   299 => x"f4c24974",
   300 => x"c481bfd5",
   301 => x"e5f4c291",
   302 => x"9a797281",
   303 => x"7287d202",
   304 => x"7189c149",
   305 => x"c1486e9a",
   306 => x"727e7080",
   307 => x"eeff059a",
   308 => x"c284c187",
   309 => x"ff04acb7",
   310 => x"486e87c9",
   311 => x"a8b7fcc0",
   312 => x"87ffc804",
   313 => x"4a744cc0",
   314 => x"c48266c4",
   315 => x"e5f4c292",
   316 => x"c8497482",
   317 => x"91c48166",
   318 => x"81e5f4c2",
   319 => x"49694a6a",
   320 => x"4b74b972",
   321 => x"bfd5f4c2",
   322 => x"c293c483",
   323 => x"6b83e5f4",
   324 => x"714872ba",
   325 => x"58a6d098",
   326 => x"f4c24974",
   327 => x"c481bfd5",
   328 => x"e5f4c291",
   329 => x"d07e6981",
   330 => x"78c048a6",
   331 => x"df4966cc",
   332 => x"c0c70229",
   333 => x"c04a7487",
   334 => x"66d092e0",
   335 => x"48ffc082",
   336 => x"4a708872",
   337 => x"c048a6d4",
   338 => x"c080c478",
   339 => x"df496e78",
   340 => x"a6e0c029",
   341 => x"d1f4c259",
   342 => x"7278c148",
   343 => x"b731c349",
   344 => x"c0b1722a",
   345 => x"91c499ff",
   346 => x"4dc5dec2",
   347 => x"4b6d8571",
   348 => x"c0c0c449",
   349 => x"f3c00299",
   350 => x"0266dc87",
   351 => x"80c887c8",
   352 => x"c57840c0",
   353 => x"f4c287ef",
   354 => x"78c148d9",
   355 => x"bfddf4c2",
   356 => x"87e1c505",
   357 => x"f81ed8c1",
   358 => x"e3f949a0",
   359 => x"1ed8c587",
   360 => x"49d1f4c2",
   361 => x"c887d9f9",
   362 => x"87c9c586",
   363 => x"d80266dc",
   364 => x"c2497387",
   365 => x"0299c0c0",
   366 => x"d087c3c0",
   367 => x"486d2bb7",
   368 => x"98fffffd",
   369 => x"fac07d70",
   370 => x"d9f4c287",
   371 => x"f2c002bf",
   372 => x"d0487387",
   373 => x"e4c028b7",
   374 => x"987058a6",
   375 => x"87e3c002",
   376 => x"bfe1f4c2",
   377 => x"c0e0c049",
   378 => x"cac00299",
   379 => x"c0497087",
   380 => x"0299c0e0",
   381 => x"6d87ccc0",
   382 => x"c0c0c248",
   383 => x"c07d70b0",
   384 => x"734b66e0",
   385 => x"c0c0c849",
   386 => x"c7c20299",
   387 => x"e1f4c287",
   388 => x"c0cc4abf",
   389 => x"cfc0029a",
   390 => x"8ac0c487",
   391 => x"87d8c002",
   392 => x"f9c0028a",
   393 => x"87ddc187",
   394 => x"ffc34973",
   395 => x"c291c299",
   396 => x"1181f9dd",
   397 => x"87dcc14b",
   398 => x"ffc34973",
   399 => x"c291c299",
   400 => x"c181f9dd",
   401 => x"dc4b1181",
   402 => x"c8c00266",
   403 => x"48a6d887",
   404 => x"ffc078d2",
   405 => x"48a6d487",
   406 => x"c078d2c4",
   407 => x"497387f6",
   408 => x"c299ffc3",
   409 => x"f9ddc291",
   410 => x"1181c181",
   411 => x"0266dc4b",
   412 => x"d887c9c0",
   413 => x"d9c148a6",
   414 => x"87d8c078",
   415 => x"c548a6d4",
   416 => x"cfc078d9",
   417 => x"c3497387",
   418 => x"91c299ff",
   419 => x"81f9ddc2",
   420 => x"4b1181c1",
   421 => x"c00266dc",
   422 => x"497387dc",
   423 => x"fcc7b9ff",
   424 => x"487199c0",
   425 => x"bfe1f4c2",
   426 => x"e5f4c298",
   427 => x"9bffc358",
   428 => x"c0b3c0c4",
   429 => x"497387d4",
   430 => x"99c0fcc7",
   431 => x"f4c24871",
   432 => x"c2b0bfe1",
   433 => x"c358e5f4",
   434 => x"66d49bff",
   435 => x"87cac002",
   436 => x"d1f4c21e",
   437 => x"87e8f449",
   438 => x"1e7386c4",
   439 => x"49d1f4c2",
   440 => x"c487ddf4",
   441 => x"0266d886",
   442 => x"1e87cac0",
   443 => x"49d1f4c2",
   444 => x"c487cdf4",
   445 => x"4866cc86",
   446 => x"a6d030c1",
   447 => x"c1486e58",
   448 => x"d07e7030",
   449 => x"80c14866",
   450 => x"c058a6d4",
   451 => x"04a8b7e0",
   452 => x"c187d9f8",
   453 => x"acb7c284",
   454 => x"87caf704",
   455 => x"48d5f4c2",
   456 => x"ff7866c4",
   457 => x"4d268edc",
   458 => x"4b264c26",
   459 => x"00004f26",
   460 => x"c01e0000",
   461 => x"c449724a",
   462 => x"e5f4c291",
   463 => x"c179ff81",
   464 => x"aab7c682",
   465 => x"c287ee04",
   466 => x"c048d5f4",
   467 => x"80c87840",
   468 => x"4f2678c0",
   469 => x"711e731e",
   470 => x"f5ddc24b",
   471 => x"87c905bf",
   472 => x"48f5ddc2",
   473 => x"c9ff78c1",
   474 => x"87dcf387",
   475 => x"c8ff4973",
   476 => x"f5fe87fc",
   477 => x"00000087",
   478 => x"f2ebf400",
   479 => x"040605f5",
   480 => x"830b030c",
   481 => x"fc00660a",
   482 => x"da005a00",
   483 => x"94800000",
   484 => x"78800508",
   485 => x"01800200",
   486 => x"09800300",
   487 => x"00800400",
   488 => x"91800100",
   489 => x"04002608",
   490 => x"00001d00",
   491 => x"00001c00",
   492 => x"0c002500",
   493 => x"00001a00",
   494 => x"00001b00",
   495 => x"00002400",
   496 => x"00011200",
   497 => x"03002e00",
   498 => x"00002d00",
   499 => x"00002300",
   500 => x"0b003600",
   501 => x"00002100",
   502 => x"00002b00",
   503 => x"00002c00",
   504 => x"00002200",
   505 => x"6c003d00",
   506 => x"00003500",
   507 => x"00003400",
   508 => x"75003e00",
   509 => x"00003200",
   510 => x"00003300",
   511 => x"6b003c00",
   512 => x"00002a00",
   513 => x"01004600",
   514 => x"73004300",
   515 => x"69003b00",
   516 => x"09004500",
   517 => x"70003a00",
   518 => x"72004200",
   519 => x"74004400",
   520 => x"00003100",
   521 => x"00005500",
   522 => x"7c004d00",
   523 => x"7a004b00",
   524 => x"00007b00",
   525 => x"71004900",
   526 => x"84004c00",
   527 => x"77005400",
   528 => x"00004100",
   529 => x"00006100",
   530 => x"7c005b00",
   531 => x"00005200",
   532 => x"0000f100",
   533 => x"00025900",
   534 => x"5d000e00",
   535 => x"00005d00",
   536 => x"79004a00",
   537 => x"05001600",
   538 => x"07007600",
   539 => x"0d000d00",
   540 => x"06001e00",
   541 => x"00002900",
   542 => x"00041400",
   543 => x"00001500",
   544 => x"00400000",
   545 => x"00400000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
