library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8f5c287",
    12 => x"86c0c84e",
    13 => x"49d8f5c2",
    14 => x"48c8e2c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dbdf",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"9a721e73",
    47 => x"87e7c002",
    48 => x"4bc148c0",
    49 => x"d106a972",
    50 => x"06827287",
    51 => x"837387c9",
    52 => x"f401a972",
    53 => x"c187c387",
    54 => x"a9723ab2",
    55 => x"80738903",
    56 => x"2b2ac107",
    57 => x"2687f305",
    58 => x"1e4f264b",
    59 => x"4dc41e75",
    60 => x"04a1b771",
    61 => x"81c1b9ff",
    62 => x"7207bdc3",
    63 => x"ff04a2b7",
    64 => x"c182c1ba",
    65 => x"eefe07bd",
    66 => x"042dc187",
    67 => x"80c1b8ff",
    68 => x"ff042d07",
    69 => x"0781c1b9",
    70 => x"4f264d26",
    71 => x"c44a711e",
    72 => x"c1484966",
    73 => x"58a6c888",
    74 => x"d6029971",
    75 => x"48d4ff87",
    76 => x"6878ffc3",
    77 => x"4966c452",
    78 => x"c888c148",
    79 => x"997158a6",
    80 => x"2687ea05",
    81 => x"1e731e4f",
    82 => x"c34bd4ff",
    83 => x"4a6b7bff",
    84 => x"6b7bffc3",
    85 => x"7232c849",
    86 => x"7bffc3b1",
    87 => x"31c84a6b",
    88 => x"ffc3b271",
    89 => x"c8496b7b",
    90 => x"71b17232",
    91 => x"2687c448",
    92 => x"264c264d",
    93 => x"0e4f264b",
    94 => x"5d5c5b5e",
    95 => x"ff4a710e",
    96 => x"49724cd4",
    97 => x"7199ffc3",
    98 => x"c8e2c27c",
    99 => x"87c805bf",
   100 => x"c94866d0",
   101 => x"58a6d430",
   102 => x"d84966d0",
   103 => x"99ffc329",
   104 => x"66d07c71",
   105 => x"c329d049",
   106 => x"7c7199ff",
   107 => x"c84966d0",
   108 => x"99ffc329",
   109 => x"66d07c71",
   110 => x"99ffc349",
   111 => x"49727c71",
   112 => x"ffc329d0",
   113 => x"6c7c7199",
   114 => x"fff0c94b",
   115 => x"abffc34d",
   116 => x"c387d005",
   117 => x"4b6c7cff",
   118 => x"c6028dc1",
   119 => x"abffc387",
   120 => x"7387f002",
   121 => x"87c7fe48",
   122 => x"ff49c01e",
   123 => x"ffc348d4",
   124 => x"c381c178",
   125 => x"04a9b7c8",
   126 => x"4f2687f1",
   127 => x"e71e731e",
   128 => x"dff8c487",
   129 => x"c01ec04b",
   130 => x"f7c1f0ff",
   131 => x"87e7fd49",
   132 => x"a8c186c4",
   133 => x"87eac005",
   134 => x"c348d4ff",
   135 => x"c0c178ff",
   136 => x"c0c0c0c0",
   137 => x"f0e1c01e",
   138 => x"fd49e9c1",
   139 => x"86c487c9",
   140 => x"ca059870",
   141 => x"48d4ff87",
   142 => x"c178ffc3",
   143 => x"fe87cb48",
   144 => x"8bc187e6",
   145 => x"87fdfe05",
   146 => x"e6fc48c0",
   147 => x"1e731e87",
   148 => x"c348d4ff",
   149 => x"4bd378ff",
   150 => x"ffc01ec0",
   151 => x"49c1c1f0",
   152 => x"c487d4fc",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187f1fd",
   158 => x"dbff058b",
   159 => x"fb48c087",
   160 => x"5e0e87f1",
   161 => x"ff0e5c5b",
   162 => x"dbfd4cd4",
   163 => x"1eeac687",
   164 => x"c1f0e1c0",
   165 => x"defb49c8",
   166 => x"c186c487",
   167 => x"87c802a8",
   168 => x"c087eafe",
   169 => x"87e2c148",
   170 => x"7087dafa",
   171 => x"ffffcf49",
   172 => x"a9eac699",
   173 => x"fe87c802",
   174 => x"48c087d3",
   175 => x"c387cbc1",
   176 => x"f1c07cff",
   177 => x"87f4fc4b",
   178 => x"c0029870",
   179 => x"1ec087eb",
   180 => x"c1f0ffc0",
   181 => x"defa49fa",
   182 => x"7086c487",
   183 => x"87d90598",
   184 => x"6c7cffc3",
   185 => x"7cffc349",
   186 => x"c17c7c7c",
   187 => x"c40299c0",
   188 => x"d548c187",
   189 => x"d148c087",
   190 => x"05abc287",
   191 => x"48c087c4",
   192 => x"8bc187c8",
   193 => x"87fdfe05",
   194 => x"e4f948c0",
   195 => x"1e731e87",
   196 => x"48c8e2c2",
   197 => x"4bc778c1",
   198 => x"c248d0ff",
   199 => x"87c8fb78",
   200 => x"c348d0ff",
   201 => x"c01ec078",
   202 => x"c0c1d0e5",
   203 => x"87c7f949",
   204 => x"a8c186c4",
   205 => x"4b87c105",
   206 => x"c505abc2",
   207 => x"c048c087",
   208 => x"8bc187f9",
   209 => x"87d0ff05",
   210 => x"c287f7fc",
   211 => x"7058cce2",
   212 => x"87cd0598",
   213 => x"ffc01ec1",
   214 => x"49d0c1f0",
   215 => x"c487d8f8",
   216 => x"48d4ff86",
   217 => x"c278ffc3",
   218 => x"e2c287fc",
   219 => x"d0ff58d0",
   220 => x"ff78c248",
   221 => x"ffc348d4",
   222 => x"f748c178",
   223 => x"5e0e87f5",
   224 => x"0e5d5c5b",
   225 => x"4cc04b71",
   226 => x"dfcdeec5",
   227 => x"48d4ff4a",
   228 => x"6878ffc3",
   229 => x"a9fec349",
   230 => x"87fdc005",
   231 => x"9b734d70",
   232 => x"d087cc02",
   233 => x"49731e66",
   234 => x"c487f1f5",
   235 => x"ff87d686",
   236 => x"d1c448d0",
   237 => x"7dffc378",
   238 => x"c14866d0",
   239 => x"58a6d488",
   240 => x"f0059870",
   241 => x"48d4ff87",
   242 => x"7878ffc3",
   243 => x"c5059b73",
   244 => x"48d0ff87",
   245 => x"4ac178d0",
   246 => x"058ac14c",
   247 => x"7487eefe",
   248 => x"87cbf648",
   249 => x"711e731e",
   250 => x"ff4bc04a",
   251 => x"ffc348d4",
   252 => x"48d0ff78",
   253 => x"ff78c3c4",
   254 => x"ffc348d4",
   255 => x"c01e7278",
   256 => x"d1c1f0ff",
   257 => x"87eff549",
   258 => x"987086c4",
   259 => x"c887d205",
   260 => x"66cc1ec0",
   261 => x"87e6fd49",
   262 => x"4b7086c4",
   263 => x"c248d0ff",
   264 => x"f5487378",
   265 => x"5e0e87cd",
   266 => x"0e5d5c5b",
   267 => x"ffc01ec0",
   268 => x"49c9c1f0",
   269 => x"d287c0f5",
   270 => x"d0e2c21e",
   271 => x"87fefc49",
   272 => x"4cc086c8",
   273 => x"b7d284c1",
   274 => x"87f804ac",
   275 => x"97d0e2c2",
   276 => x"c0c349bf",
   277 => x"a9c0c199",
   278 => x"87e7c005",
   279 => x"97d7e2c2",
   280 => x"31d049bf",
   281 => x"97d8e2c2",
   282 => x"32c84abf",
   283 => x"e2c2b172",
   284 => x"4abf97d9",
   285 => x"cf4c71b1",
   286 => x"9cffffff",
   287 => x"34ca84c1",
   288 => x"c287e7c1",
   289 => x"bf97d9e2",
   290 => x"c631c149",
   291 => x"dae2c299",
   292 => x"c74abf97",
   293 => x"b1722ab7",
   294 => x"97d5e2c2",
   295 => x"cf4d4abf",
   296 => x"d6e2c29d",
   297 => x"c34abf97",
   298 => x"c232ca9a",
   299 => x"bf97d7e2",
   300 => x"7333c24b",
   301 => x"d8e2c2b2",
   302 => x"c34bbf97",
   303 => x"b7c69bc0",
   304 => x"c2b2732b",
   305 => x"7148c181",
   306 => x"c1497030",
   307 => x"70307548",
   308 => x"c14c724d",
   309 => x"c8947184",
   310 => x"06adb7c0",
   311 => x"34c187cc",
   312 => x"c0c82db7",
   313 => x"ff01adb7",
   314 => x"487487f4",
   315 => x"0e87c0f2",
   316 => x"5d5c5b5e",
   317 => x"c286f80e",
   318 => x"c048f6ea",
   319 => x"eee2c278",
   320 => x"fb49c01e",
   321 => x"86c487de",
   322 => x"c5059870",
   323 => x"c948c087",
   324 => x"4dc087ce",
   325 => x"efc07ec1",
   326 => x"c249bfd8",
   327 => x"714ae4e3",
   328 => x"c4ed4bc8",
   329 => x"05987087",
   330 => x"7ec087c2",
   331 => x"bfd4efc0",
   332 => x"c0e4c249",
   333 => x"4bc8714a",
   334 => x"7087eeec",
   335 => x"87c20598",
   336 => x"026e7ec0",
   337 => x"c287fdc0",
   338 => x"4dbff4e9",
   339 => x"9feceac2",
   340 => x"c5487ebf",
   341 => x"05a8ead6",
   342 => x"e9c287c7",
   343 => x"ce4dbff4",
   344 => x"ca486e87",
   345 => x"02a8d5e9",
   346 => x"48c087c5",
   347 => x"c287f1c7",
   348 => x"751eeee2",
   349 => x"87ecf949",
   350 => x"987086c4",
   351 => x"c087c505",
   352 => x"87dcc748",
   353 => x"bfd4efc0",
   354 => x"c0e4c249",
   355 => x"4bc8714a",
   356 => x"7087d6eb",
   357 => x"87c80598",
   358 => x"48f6eac2",
   359 => x"87da78c1",
   360 => x"bfd8efc0",
   361 => x"e4e3c249",
   362 => x"4bc8714a",
   363 => x"7087faea",
   364 => x"c5c00298",
   365 => x"c648c087",
   366 => x"eac287e6",
   367 => x"49bf97ec",
   368 => x"05a9d5c1",
   369 => x"c287cdc0",
   370 => x"bf97edea",
   371 => x"a9eac249",
   372 => x"87c5c002",
   373 => x"c7c648c0",
   374 => x"eee2c287",
   375 => x"487ebf97",
   376 => x"02a8e9c3",
   377 => x"6e87cec0",
   378 => x"a8ebc348",
   379 => x"87c5c002",
   380 => x"ebc548c0",
   381 => x"f9e2c287",
   382 => x"9949bf97",
   383 => x"87ccc005",
   384 => x"97fae2c2",
   385 => x"a9c249bf",
   386 => x"87c5c002",
   387 => x"cfc548c0",
   388 => x"fbe2c287",
   389 => x"c248bf97",
   390 => x"7058f2ea",
   391 => x"88c1484c",
   392 => x"58f6eac2",
   393 => x"97fce2c2",
   394 => x"817549bf",
   395 => x"97fde2c2",
   396 => x"32c84abf",
   397 => x"c27ea172",
   398 => x"6e48c3ef",
   399 => x"fee2c278",
   400 => x"c848bf97",
   401 => x"eac258a6",
   402 => x"c202bff6",
   403 => x"efc087d4",
   404 => x"c249bfd4",
   405 => x"714ac0e4",
   406 => x"cce84bc8",
   407 => x"02987087",
   408 => x"c087c5c0",
   409 => x"87f8c348",
   410 => x"bfeeeac2",
   411 => x"d7efc24c",
   412 => x"d3e3c25c",
   413 => x"c849bf97",
   414 => x"d2e3c231",
   415 => x"a14abf97",
   416 => x"d4e3c249",
   417 => x"d04abf97",
   418 => x"49a17232",
   419 => x"97d5e3c2",
   420 => x"32d84abf",
   421 => x"c449a172",
   422 => x"efc29166",
   423 => x"c281bfc3",
   424 => x"c259cbef",
   425 => x"bf97dbe3",
   426 => x"c232c84a",
   427 => x"bf97dae3",
   428 => x"c24aa24b",
   429 => x"bf97dce3",
   430 => x"7333d04b",
   431 => x"e3c24aa2",
   432 => x"4bbf97dd",
   433 => x"33d89bcf",
   434 => x"c24aa273",
   435 => x"c25acfef",
   436 => x"4abfcbef",
   437 => x"92748ac2",
   438 => x"48cfefc2",
   439 => x"c178a172",
   440 => x"e3c287ca",
   441 => x"49bf97c0",
   442 => x"e2c231c8",
   443 => x"4abf97ff",
   444 => x"eac249a1",
   445 => x"eac259fe",
   446 => x"c549bffa",
   447 => x"81ffc731",
   448 => x"efc229c9",
   449 => x"e3c259d7",
   450 => x"4abf97c5",
   451 => x"e3c232c8",
   452 => x"4bbf97c4",
   453 => x"66c44aa2",
   454 => x"c2826e92",
   455 => x"c25ad3ef",
   456 => x"c048cbef",
   457 => x"c7efc278",
   458 => x"78a17248",
   459 => x"48d7efc2",
   460 => x"bfcbefc2",
   461 => x"dbefc278",
   462 => x"cfefc248",
   463 => x"eac278bf",
   464 => x"c002bff6",
   465 => x"487487c9",
   466 => x"7e7030c4",
   467 => x"c287c9c0",
   468 => x"48bfd3ef",
   469 => x"7e7030c4",
   470 => x"48faeac2",
   471 => x"48c1786e",
   472 => x"4d268ef8",
   473 => x"4b264c26",
   474 => x"5e0e4f26",
   475 => x"0e5d5c5b",
   476 => x"eac24a71",
   477 => x"cb02bff6",
   478 => x"c74b7287",
   479 => x"c14c722b",
   480 => x"87c99cff",
   481 => x"2bc84b72",
   482 => x"ffc34c72",
   483 => x"c3efc29c",
   484 => x"efc083bf",
   485 => x"02abbfd0",
   486 => x"efc087d9",
   487 => x"e2c25bd4",
   488 => x"49731eee",
   489 => x"c487fdf0",
   490 => x"05987086",
   491 => x"48c087c5",
   492 => x"c287e6c0",
   493 => x"02bff6ea",
   494 => x"497487d2",
   495 => x"e2c291c4",
   496 => x"4d6981ee",
   497 => x"ffffffcf",
   498 => x"87cb9dff",
   499 => x"91c24974",
   500 => x"81eee2c2",
   501 => x"754d699f",
   502 => x"87c6fe48",
   503 => x"5c5b5e0e",
   504 => x"86f80e5d",
   505 => x"059c4c71",
   506 => x"48c087c5",
   507 => x"c887c2c3",
   508 => x"486e7ea4",
   509 => x"66d878c0",
   510 => x"d887c702",
   511 => x"05bf9766",
   512 => x"48c087c5",
   513 => x"c087eac2",
   514 => x"4949c11e",
   515 => x"c487e6c7",
   516 => x"9d4d7086",
   517 => x"87c2c102",
   518 => x"4afeeac2",
   519 => x"e04966d8",
   520 => x"987087ec",
   521 => x"87f2c002",
   522 => x"66d84a75",
   523 => x"e14bcb49",
   524 => x"987087d1",
   525 => x"87e2c002",
   526 => x"9d751ec0",
   527 => x"c887c702",
   528 => x"78c048a6",
   529 => x"a6c887c5",
   530 => x"c878c148",
   531 => x"e4c64966",
   532 => x"7086c487",
   533 => x"fe059d4d",
   534 => x"9d7587fe",
   535 => x"87cfc102",
   536 => x"6e49a5dc",
   537 => x"da786948",
   538 => x"a6c449a5",
   539 => x"78a4c448",
   540 => x"c448699f",
   541 => x"c2780866",
   542 => x"02bff6ea",
   543 => x"a5d487d2",
   544 => x"49699f49",
   545 => x"99ffffc0",
   546 => x"30d04871",
   547 => x"87c27e70",
   548 => x"496e7ec0",
   549 => x"bf66c448",
   550 => x"0866c480",
   551 => x"cc7cc078",
   552 => x"66c449a4",
   553 => x"a4d079bf",
   554 => x"c179c049",
   555 => x"c087c248",
   556 => x"fa8ef848",
   557 => x"5e0e87ec",
   558 => x"0e5d5c5b",
   559 => x"029c4c71",
   560 => x"c887cac1",
   561 => x"026949a4",
   562 => x"d087c2c1",
   563 => x"496c4a66",
   564 => x"5aa6d482",
   565 => x"b94d66d0",
   566 => x"bff2eac2",
   567 => x"72baff4a",
   568 => x"02997199",
   569 => x"c487e4c0",
   570 => x"496b4ba4",
   571 => x"7087fbf9",
   572 => x"eeeac27b",
   573 => x"816c49bf",
   574 => x"b9757c71",
   575 => x"bff2eac2",
   576 => x"72baff4a",
   577 => x"05997199",
   578 => x"7587dcff",
   579 => x"87d2f97c",
   580 => x"711e731e",
   581 => x"c7029b4b",
   582 => x"49a3c887",
   583 => x"87c50569",
   584 => x"f7c048c0",
   585 => x"c7efc287",
   586 => x"a3c44abf",
   587 => x"c2496949",
   588 => x"eeeac289",
   589 => x"a27191bf",
   590 => x"f2eac24a",
   591 => x"996b49bf",
   592 => x"c04aa271",
   593 => x"c85ad4ef",
   594 => x"49721e66",
   595 => x"c487d5ea",
   596 => x"05987086",
   597 => x"48c087c4",
   598 => x"48c187c2",
   599 => x"1e87c7f8",
   600 => x"4b711e73",
   601 => x"e4c0029b",
   602 => x"dbefc287",
   603 => x"c24a735b",
   604 => x"eeeac28a",
   605 => x"c29249bf",
   606 => x"48bfc7ef",
   607 => x"efc28072",
   608 => x"487158df",
   609 => x"eac230c4",
   610 => x"edc058fe",
   611 => x"d7efc287",
   612 => x"cbefc248",
   613 => x"efc278bf",
   614 => x"efc248db",
   615 => x"c278bfcf",
   616 => x"02bff6ea",
   617 => x"eac287c9",
   618 => x"c449bfee",
   619 => x"c287c731",
   620 => x"49bfd3ef",
   621 => x"eac231c4",
   622 => x"e9f659fe",
   623 => x"5b5e0e87",
   624 => x"4a710e5c",
   625 => x"9a724bc0",
   626 => x"87e1c002",
   627 => x"9f49a2da",
   628 => x"eac24b69",
   629 => x"cf02bff6",
   630 => x"49a2d487",
   631 => x"4c49699f",
   632 => x"9cffffc0",
   633 => x"87c234d0",
   634 => x"49744cc0",
   635 => x"fd4973b3",
   636 => x"eff587ed",
   637 => x"5b5e0e87",
   638 => x"f40e5d5c",
   639 => x"c04a7186",
   640 => x"029a727e",
   641 => x"e2c287d8",
   642 => x"78c048ea",
   643 => x"48e2e2c2",
   644 => x"bfdbefc2",
   645 => x"e6e2c278",
   646 => x"d7efc248",
   647 => x"ebc278bf",
   648 => x"50c048cb",
   649 => x"bffaeac2",
   650 => x"eae2c249",
   651 => x"aa714abf",
   652 => x"87c9c403",
   653 => x"99cf4972",
   654 => x"87e9c005",
   655 => x"48d0efc0",
   656 => x"bfe2e2c2",
   657 => x"eee2c278",
   658 => x"e2e2c21e",
   659 => x"e2c249bf",
   660 => x"a1c148e2",
   661 => x"cbe67178",
   662 => x"c086c487",
   663 => x"c248ccef",
   664 => x"cc78eee2",
   665 => x"ccefc087",
   666 => x"e0c048bf",
   667 => x"d0efc080",
   668 => x"eae2c258",
   669 => x"80c148bf",
   670 => x"58eee2c2",
   671 => x"000bcc27",
   672 => x"bf97bf00",
   673 => x"c2029d4d",
   674 => x"e5c387e3",
   675 => x"dcc202ad",
   676 => x"ccefc087",
   677 => x"a3cb4bbf",
   678 => x"cf4c1149",
   679 => x"d2c105ac",
   680 => x"df497587",
   681 => x"cd89c199",
   682 => x"feeac291",
   683 => x"4aa3c181",
   684 => x"a3c35112",
   685 => x"c551124a",
   686 => x"51124aa3",
   687 => x"124aa3c7",
   688 => x"4aa3c951",
   689 => x"a3ce5112",
   690 => x"d051124a",
   691 => x"51124aa3",
   692 => x"124aa3d2",
   693 => x"4aa3d451",
   694 => x"a3d65112",
   695 => x"d851124a",
   696 => x"51124aa3",
   697 => x"124aa3dc",
   698 => x"4aa3de51",
   699 => x"7ec15112",
   700 => x"7487fac0",
   701 => x"0599c849",
   702 => x"7487ebc0",
   703 => x"0599d049",
   704 => x"66dc87d1",
   705 => x"87cbc002",
   706 => x"66dc4973",
   707 => x"0298700f",
   708 => x"6e87d3c0",
   709 => x"87c6c005",
   710 => x"48feeac2",
   711 => x"efc050c0",
   712 => x"c248bfcc",
   713 => x"ebc287e1",
   714 => x"50c048cb",
   715 => x"faeac27e",
   716 => x"e2c249bf",
   717 => x"714abfea",
   718 => x"f7fb04aa",
   719 => x"dbefc287",
   720 => x"c8c005bf",
   721 => x"f6eac287",
   722 => x"f8c102bf",
   723 => x"e6e2c287",
   724 => x"d5f049bf",
   725 => x"c2497087",
   726 => x"c459eae2",
   727 => x"e2c248a6",
   728 => x"c278bfe6",
   729 => x"02bff6ea",
   730 => x"c487d8c0",
   731 => x"ffcf4966",
   732 => x"99f8ffff",
   733 => x"c5c002a9",
   734 => x"c04cc087",
   735 => x"4cc187e1",
   736 => x"c487dcc0",
   737 => x"ffcf4966",
   738 => x"02a999f8",
   739 => x"c887c8c0",
   740 => x"78c048a6",
   741 => x"c887c5c0",
   742 => x"78c148a6",
   743 => x"744c66c8",
   744 => x"e0c0059c",
   745 => x"4966c487",
   746 => x"eac289c2",
   747 => x"914abfee",
   748 => x"bfc7efc2",
   749 => x"e2e2c24a",
   750 => x"78a17248",
   751 => x"48eae2c2",
   752 => x"dff978c0",
   753 => x"f448c087",
   754 => x"87d6ee8e",
   755 => x"00000000",
   756 => x"ffffffff",
   757 => x"00000bdc",
   758 => x"00000be5",
   759 => x"33544146",
   760 => x"20202032",
   761 => x"54414600",
   762 => x"20203631",
   763 => x"ff1e0020",
   764 => x"ffc348d4",
   765 => x"26486878",
   766 => x"d4ff1e4f",
   767 => x"78ffc348",
   768 => x"c048d0ff",
   769 => x"d4ff78e1",
   770 => x"c278d448",
   771 => x"ff48dfef",
   772 => x"2650bfd4",
   773 => x"d0ff1e4f",
   774 => x"78e0c048",
   775 => x"ff1e4f26",
   776 => x"497087cc",
   777 => x"87c60299",
   778 => x"05a9fbc0",
   779 => x"487187f1",
   780 => x"5e0e4f26",
   781 => x"710e5c5b",
   782 => x"fe4cc04b",
   783 => x"497087f0",
   784 => x"f9c00299",
   785 => x"a9ecc087",
   786 => x"87f2c002",
   787 => x"02a9fbc0",
   788 => x"cc87ebc0",
   789 => x"03acb766",
   790 => x"66d087c7",
   791 => x"7187c202",
   792 => x"02997153",
   793 => x"84c187c2",
   794 => x"7087c3fe",
   795 => x"cd029949",
   796 => x"a9ecc087",
   797 => x"c087c702",
   798 => x"ff05a9fb",
   799 => x"66d087d5",
   800 => x"c087c302",
   801 => x"ecc07b97",
   802 => x"87c405a9",
   803 => x"87c54a74",
   804 => x"0ac04a74",
   805 => x"c248728a",
   806 => x"264d2687",
   807 => x"264b264c",
   808 => x"c9fd1e4f",
   809 => x"4a497087",
   810 => x"04aaf0c0",
   811 => x"f9c087c9",
   812 => x"87c301aa",
   813 => x"c18af0c0",
   814 => x"c904aac1",
   815 => x"aadac187",
   816 => x"c087c301",
   817 => x"48728af7",
   818 => x"5e0e4f26",
   819 => x"710e5c5b",
   820 => x"4bd4ff4a",
   821 => x"e7c04972",
   822 => x"9c4c7087",
   823 => x"c187c202",
   824 => x"48d0ff8c",
   825 => x"d5c178c5",
   826 => x"c649747b",
   827 => x"fce0c131",
   828 => x"484abf97",
   829 => x"7b70b071",
   830 => x"c448d0ff",
   831 => x"87dbfe78",
   832 => x"5c5b5e0e",
   833 => x"86f80e5d",
   834 => x"7ec04c71",
   835 => x"c087eafb",
   836 => x"edf6c04b",
   837 => x"c049bf97",
   838 => x"87cf04a9",
   839 => x"c187fffb",
   840 => x"edf6c083",
   841 => x"ab49bf97",
   842 => x"c087f106",
   843 => x"bf97edf6",
   844 => x"fa87cf02",
   845 => x"497087f8",
   846 => x"87c60299",
   847 => x"05a9ecc0",
   848 => x"4bc087f1",
   849 => x"7087e7fa",
   850 => x"87e2fa4d",
   851 => x"fa58a6c8",
   852 => x"4a7087dc",
   853 => x"a4c883c1",
   854 => x"49699749",
   855 => x"87c702ad",
   856 => x"05adffc0",
   857 => x"c987e7c0",
   858 => x"699749a4",
   859 => x"a966c449",
   860 => x"4887c702",
   861 => x"05a8ffc0",
   862 => x"a4ca87d4",
   863 => x"49699749",
   864 => x"87c602aa",
   865 => x"05aaffc0",
   866 => x"7ec187c4",
   867 => x"ecc087d0",
   868 => x"87c602ad",
   869 => x"05adfbc0",
   870 => x"4bc087c4",
   871 => x"026e7ec1",
   872 => x"f987e1fe",
   873 => x"487387ef",
   874 => x"ecfb8ef8",
   875 => x"5e0e0087",
   876 => x"0e5d5c5b",
   877 => x"4d7186f8",
   878 => x"754bd4ff",
   879 => x"e4efc21e",
   880 => x"87d8e849",
   881 => x"987086c4",
   882 => x"87ccc402",
   883 => x"c148a6c4",
   884 => x"78bffee0",
   885 => x"f1fb4975",
   886 => x"48d0ff87",
   887 => x"d6c178c5",
   888 => x"754ac07b",
   889 => x"7b1149a2",
   890 => x"b7cb82c1",
   891 => x"87f304aa",
   892 => x"ffc34acc",
   893 => x"c082c17b",
   894 => x"04aab7e0",
   895 => x"d0ff87f4",
   896 => x"c378c448",
   897 => x"78c57bff",
   898 => x"c17bd3c1",
   899 => x"6678c47b",
   900 => x"a8b7c048",
   901 => x"87f0c206",
   902 => x"bfecefc2",
   903 => x"4866c44c",
   904 => x"a6c88874",
   905 => x"029c7458",
   906 => x"c287f9c1",
   907 => x"c87eeee2",
   908 => x"c08c4dc0",
   909 => x"c603acb7",
   910 => x"a4c0c887",
   911 => x"c24cc04d",
   912 => x"bf97dfef",
   913 => x"0299d049",
   914 => x"1ec087d1",
   915 => x"49e4efc2",
   916 => x"c487fdea",
   917 => x"4a497086",
   918 => x"c287eec0",
   919 => x"c21eeee2",
   920 => x"ea49e4ef",
   921 => x"86c487ea",
   922 => x"ff4a4970",
   923 => x"c5c848d0",
   924 => x"7bd4c178",
   925 => x"7bbf976e",
   926 => x"80c1486e",
   927 => x"8dc17e70",
   928 => x"87f0ff05",
   929 => x"c448d0ff",
   930 => x"059a7278",
   931 => x"48c087c5",
   932 => x"c187c7c1",
   933 => x"e4efc21e",
   934 => x"87dae849",
   935 => x"9c7486c4",
   936 => x"87c7fe05",
   937 => x"c04866c4",
   938 => x"d106a8b7",
   939 => x"e4efc287",
   940 => x"d078c048",
   941 => x"f478c080",
   942 => x"f0efc280",
   943 => x"66c478bf",
   944 => x"a8b7c048",
   945 => x"87d0fd01",
   946 => x"c548d0ff",
   947 => x"7bd3c178",
   948 => x"78c47bc0",
   949 => x"87c248c1",
   950 => x"8ef848c0",
   951 => x"4c264d26",
   952 => x"4f264b26",
   953 => x"5c5b5e0e",
   954 => x"711e0e5d",
   955 => x"4d4cc04b",
   956 => x"e8c004ab",
   957 => x"c0f4c087",
   958 => x"029d751e",
   959 => x"4ac087c4",
   960 => x"4ac187c2",
   961 => x"eceb4972",
   962 => x"7086c487",
   963 => x"6e84c17e",
   964 => x"7387c205",
   965 => x"7385c14c",
   966 => x"d8ff06ac",
   967 => x"26486e87",
   968 => x"1e87f9fe",
   969 => x"66c44a71",
   970 => x"7287c505",
   971 => x"87fef949",
   972 => x"5e0e4f26",
   973 => x"0e5d5c5b",
   974 => x"494c711e",
   975 => x"f0c291de",
   976 => x"85714dcc",
   977 => x"c1026d97",
   978 => x"efc287dd",
   979 => x"744abff8",
   980 => x"fe497282",
   981 => x"7e7087ce",
   982 => x"c0029848",
   983 => x"f0c287f2",
   984 => x"4a704bc0",
   985 => x"c4ff49cb",
   986 => x"4b7487fd",
   987 => x"e1c193cb",
   988 => x"83c483d0",
   989 => x"7bebfec0",
   990 => x"c1c14974",
   991 => x"7b7587f3",
   992 => x"97fde0c1",
   993 => x"c21e49bf",
   994 => x"fe49c0f0",
   995 => x"86c487d5",
   996 => x"c1c14974",
   997 => x"49c087db",
   998 => x"87fac2c1",
   999 => x"48e0efc2",
  1000 => x"49c178c0",
  1001 => x"2687dcde",
  1002 => x"4c87f1fc",
  1003 => x"6964616f",
  1004 => x"2e2e676e",
  1005 => x"5e0e002e",
  1006 => x"710e5c5b",
  1007 => x"efc24a4b",
  1008 => x"7282bff8",
  1009 => x"87dcfc49",
  1010 => x"029c4c70",
  1011 => x"e74987c4",
  1012 => x"efc287eb",
  1013 => x"78c048f8",
  1014 => x"e6dd49c1",
  1015 => x"87fefb87",
  1016 => x"5c5b5e0e",
  1017 => x"86f40e5d",
  1018 => x"4deee2c2",
  1019 => x"a6c44cc0",
  1020 => x"c278c048",
  1021 => x"49bff8ef",
  1022 => x"c106a9c0",
  1023 => x"e2c287c1",
  1024 => x"029848ee",
  1025 => x"c087f8c0",
  1026 => x"c81ec0f4",
  1027 => x"87c70266",
  1028 => x"c048a6c4",
  1029 => x"c487c578",
  1030 => x"78c148a6",
  1031 => x"e74966c4",
  1032 => x"86c487d3",
  1033 => x"84c14d70",
  1034 => x"c14866c4",
  1035 => x"58a6c880",
  1036 => x"bff8efc2",
  1037 => x"c603ac49",
  1038 => x"059d7587",
  1039 => x"c087c8ff",
  1040 => x"029d754c",
  1041 => x"c087e0c3",
  1042 => x"c81ec0f4",
  1043 => x"87c70266",
  1044 => x"c048a6cc",
  1045 => x"cc87c578",
  1046 => x"78c148a6",
  1047 => x"e64966cc",
  1048 => x"86c487d3",
  1049 => x"98487e70",
  1050 => x"87e8c202",
  1051 => x"9781cb49",
  1052 => x"99d04969",
  1053 => x"87d6c102",
  1054 => x"4af6fec0",
  1055 => x"91cb4974",
  1056 => x"81d0e1c1",
  1057 => x"81c87972",
  1058 => x"7451ffc3",
  1059 => x"c291de49",
  1060 => x"714dccf0",
  1061 => x"97c1c285",
  1062 => x"49a5c17d",
  1063 => x"c251e0c0",
  1064 => x"bf97feea",
  1065 => x"c187d202",
  1066 => x"4ba5c284",
  1067 => x"4afeeac2",
  1068 => x"fffe49db",
  1069 => x"dbc187f1",
  1070 => x"49a5cd87",
  1071 => x"84c151c0",
  1072 => x"6e4ba5c2",
  1073 => x"fe49cb4a",
  1074 => x"c187dcff",
  1075 => x"fcc087c6",
  1076 => x"49744af2",
  1077 => x"e1c191cb",
  1078 => x"797281d0",
  1079 => x"97feeac2",
  1080 => x"87d802bf",
  1081 => x"91de4974",
  1082 => x"f0c284c1",
  1083 => x"83714bcc",
  1084 => x"4afeeac2",
  1085 => x"fefe49dd",
  1086 => x"87d887ed",
  1087 => x"93de4b74",
  1088 => x"83ccf0c2",
  1089 => x"c049a3cb",
  1090 => x"7384c151",
  1091 => x"49cb4a6e",
  1092 => x"87d3fefe",
  1093 => x"c14866c4",
  1094 => x"58a6c880",
  1095 => x"c003acc7",
  1096 => x"056e87c5",
  1097 => x"7487e0fc",
  1098 => x"f68ef448",
  1099 => x"731e87ee",
  1100 => x"494b711e",
  1101 => x"e1c191cb",
  1102 => x"a1c881d0",
  1103 => x"fce0c14a",
  1104 => x"c9501248",
  1105 => x"f6c04aa1",
  1106 => x"501248ed",
  1107 => x"e0c181ca",
  1108 => x"501148fd",
  1109 => x"97fde0c1",
  1110 => x"c01e49bf",
  1111 => x"87c3f749",
  1112 => x"48e0efc2",
  1113 => x"49c178de",
  1114 => x"2687d8d7",
  1115 => x"1e87f1f5",
  1116 => x"cb494a71",
  1117 => x"d0e1c191",
  1118 => x"1181c881",
  1119 => x"e4efc248",
  1120 => x"f8efc258",
  1121 => x"c178c048",
  1122 => x"87f7d649",
  1123 => x"c01e4f26",
  1124 => x"c1fbc049",
  1125 => x"1e4f2687",
  1126 => x"d2029971",
  1127 => x"e5e2c187",
  1128 => x"f750c048",
  1129 => x"efc5c180",
  1130 => x"c9e1c140",
  1131 => x"c187ce78",
  1132 => x"c148e1e2",
  1133 => x"fc78c2e1",
  1134 => x"cec6c180",
  1135 => x"0e4f2678",
  1136 => x"5d5c5b5e",
  1137 => x"7186f40e",
  1138 => x"91cb494d",
  1139 => x"81d0e1c1",
  1140 => x"ca4aa1c8",
  1141 => x"a6c47ea1",
  1142 => x"e8f3c248",
  1143 => x"976e78bf",
  1144 => x"66c44bbf",
  1145 => x"70287348",
  1146 => x"48124c4b",
  1147 => x"7058a6cc",
  1148 => x"c984c19c",
  1149 => x"49699781",
  1150 => x"c204acb7",
  1151 => x"6e4cc087",
  1152 => x"c84abf97",
  1153 => x"31724966",
  1154 => x"66c4b9ff",
  1155 => x"72487499",
  1156 => x"484a7030",
  1157 => x"f3c2b071",
  1158 => x"e5c058ec",
  1159 => x"49c087d3",
  1160 => x"7587e0d4",
  1161 => x"c8f7c049",
  1162 => x"f28ef487",
  1163 => x"731e87ee",
  1164 => x"494b711e",
  1165 => x"7387c8fe",
  1166 => x"87c3fe49",
  1167 => x"1e87e1f2",
  1168 => x"4b711e73",
  1169 => x"024aa3c6",
  1170 => x"8ac187db",
  1171 => x"8a87d602",
  1172 => x"87dac102",
  1173 => x"fcc0028a",
  1174 => x"c0028a87",
  1175 => x"028a87e1",
  1176 => x"dbc187cb",
  1177 => x"fc49c787",
  1178 => x"dec187c5",
  1179 => x"f8efc287",
  1180 => x"cbc102bf",
  1181 => x"88c14887",
  1182 => x"58fcefc2",
  1183 => x"c287c1c1",
  1184 => x"02bffcef",
  1185 => x"c287f9c0",
  1186 => x"48bff8ef",
  1187 => x"efc280c1",
  1188 => x"ebc058fc",
  1189 => x"f8efc287",
  1190 => x"89c649bf",
  1191 => x"59fcefc2",
  1192 => x"03a9b7c0",
  1193 => x"efc287da",
  1194 => x"78c048f8",
  1195 => x"efc287d2",
  1196 => x"cb02bffc",
  1197 => x"f8efc287",
  1198 => x"80c648bf",
  1199 => x"58fcefc2",
  1200 => x"fed149c0",
  1201 => x"c0497387",
  1202 => x"f087e6f4",
  1203 => x"5e0e87d2",
  1204 => x"0e5d5c5b",
  1205 => x"dc86d0ff",
  1206 => x"a6c859a6",
  1207 => x"c478c048",
  1208 => x"66c4c180",
  1209 => x"c180c478",
  1210 => x"c180c478",
  1211 => x"fcefc278",
  1212 => x"c278c148",
  1213 => x"48bfe0ef",
  1214 => x"cb05a8de",
  1215 => x"87e0f387",
  1216 => x"a6cc4970",
  1217 => x"87facf59",
  1218 => x"e487eee3",
  1219 => x"dde387d0",
  1220 => x"c04c7087",
  1221 => x"c102acfb",
  1222 => x"66d887fb",
  1223 => x"87edc105",
  1224 => x"4a66c0c1",
  1225 => x"7e6a82c4",
  1226 => x"dcc11e72",
  1227 => x"66c448f7",
  1228 => x"4aa1c849",
  1229 => x"aa714120",
  1230 => x"1087f905",
  1231 => x"c14a2651",
  1232 => x"c14866c0",
  1233 => x"6a78eec4",
  1234 => x"7481c749",
  1235 => x"66c0c151",
  1236 => x"c181c849",
  1237 => x"66c0c151",
  1238 => x"c081c949",
  1239 => x"66c0c151",
  1240 => x"c081ca49",
  1241 => x"d81ec151",
  1242 => x"c8496a1e",
  1243 => x"87c2e381",
  1244 => x"c4c186c8",
  1245 => x"a8c04866",
  1246 => x"c887c701",
  1247 => x"78c148a6",
  1248 => x"c4c187ce",
  1249 => x"88c14866",
  1250 => x"c358a6d0",
  1251 => x"87cee287",
  1252 => x"c248a6d0",
  1253 => x"029c7478",
  1254 => x"c887e3cd",
  1255 => x"c8c14866",
  1256 => x"cd03a866",
  1257 => x"a6dc87d8",
  1258 => x"e878c048",
  1259 => x"e078c080",
  1260 => x"4c7087fc",
  1261 => x"05acd0c1",
  1262 => x"c487d8c2",
  1263 => x"e0e37e66",
  1264 => x"c8497087",
  1265 => x"e5e059a6",
  1266 => x"c04c7087",
  1267 => x"c105acec",
  1268 => x"66c887ec",
  1269 => x"c191cb49",
  1270 => x"c48166c0",
  1271 => x"4d6a4aa1",
  1272 => x"c44aa1c8",
  1273 => x"c5c15266",
  1274 => x"c1e079ef",
  1275 => x"9c4c7087",
  1276 => x"c087d902",
  1277 => x"d302acfb",
  1278 => x"ff557487",
  1279 => x"7087efdf",
  1280 => x"c7029c4c",
  1281 => x"acfbc087",
  1282 => x"87edff05",
  1283 => x"c255e0c0",
  1284 => x"97c055c1",
  1285 => x"4966d87d",
  1286 => x"db05a96e",
  1287 => x"4866c887",
  1288 => x"04a866cc",
  1289 => x"66c887ca",
  1290 => x"cc80c148",
  1291 => x"87c858a6",
  1292 => x"c14866cc",
  1293 => x"58a6d088",
  1294 => x"87f2deff",
  1295 => x"d0c14c70",
  1296 => x"87c805ac",
  1297 => x"c14866d4",
  1298 => x"58a6d880",
  1299 => x"02acd0c1",
  1300 => x"c087e8fd",
  1301 => x"d848a6e0",
  1302 => x"66c47866",
  1303 => x"66e0c048",
  1304 => x"ebc905a8",
  1305 => x"a6e4c087",
  1306 => x"7478c048",
  1307 => x"88fbc048",
  1308 => x"98487e70",
  1309 => x"87edc902",
  1310 => x"7088cb48",
  1311 => x"0298487e",
  1312 => x"4887cdc1",
  1313 => x"7e7088c9",
  1314 => x"c4029848",
  1315 => x"c44887c1",
  1316 => x"487e7088",
  1317 => x"87ce0298",
  1318 => x"7088c148",
  1319 => x"0298487e",
  1320 => x"c887ecc3",
  1321 => x"a6dc87e1",
  1322 => x"78f0c048",
  1323 => x"87fedcff",
  1324 => x"ecc04c70",
  1325 => x"c4c002ac",
  1326 => x"a6e0c087",
  1327 => x"acecc05c",
  1328 => x"ff87cd02",
  1329 => x"7087e7dc",
  1330 => x"acecc04c",
  1331 => x"87f3ff05",
  1332 => x"02acecc0",
  1333 => x"ff87c4c0",
  1334 => x"c087d3dc",
  1335 => x"d01eca1e",
  1336 => x"91cb4966",
  1337 => x"4866c8c1",
  1338 => x"a6cc8071",
  1339 => x"4866c858",
  1340 => x"a6d080c4",
  1341 => x"bf66cc58",
  1342 => x"f5dcff49",
  1343 => x"de1ec187",
  1344 => x"bf66d41e",
  1345 => x"e9dcff49",
  1346 => x"7086d087",
  1347 => x"8909c049",
  1348 => x"59a6ecc0",
  1349 => x"4866e8c0",
  1350 => x"c006a8c0",
  1351 => x"e8c087ee",
  1352 => x"a8dd4866",
  1353 => x"87e4c003",
  1354 => x"49bf66c4",
  1355 => x"8166e8c0",
  1356 => x"c051e0c0",
  1357 => x"c14966e8",
  1358 => x"bf66c481",
  1359 => x"51c1c281",
  1360 => x"4966e8c0",
  1361 => x"66c481c2",
  1362 => x"51c081bf",
  1363 => x"c4c1486e",
  1364 => x"496e78ee",
  1365 => x"66d081c8",
  1366 => x"c9496e51",
  1367 => x"5166d481",
  1368 => x"81ca496e",
  1369 => x"d05166dc",
  1370 => x"80c14866",
  1371 => x"c858a6d4",
  1372 => x"66cc4866",
  1373 => x"cbc004a8",
  1374 => x"4866c887",
  1375 => x"a6cc80c1",
  1376 => x"87e1c558",
  1377 => x"c14866cc",
  1378 => x"58a6d088",
  1379 => x"ff87d6c5",
  1380 => x"7087cedc",
  1381 => x"a6ecc049",
  1382 => x"c4dcff59",
  1383 => x"c0497087",
  1384 => x"dc59a6e0",
  1385 => x"ecc04866",
  1386 => x"cac005a8",
  1387 => x"48a6dc87",
  1388 => x"7866e8c0",
  1389 => x"ff87c4c0",
  1390 => x"c887f3d8",
  1391 => x"91cb4966",
  1392 => x"4866c0c1",
  1393 => x"7e708071",
  1394 => x"6e82c84a",
  1395 => x"c081ca49",
  1396 => x"dc5166e8",
  1397 => x"81c14966",
  1398 => x"8966e8c0",
  1399 => x"307148c1",
  1400 => x"89c14970",
  1401 => x"c27a9771",
  1402 => x"49bfe8f3",
  1403 => x"2966e8c0",
  1404 => x"484a6a97",
  1405 => x"f0c09871",
  1406 => x"496e58a6",
  1407 => x"4d6981c4",
  1408 => x"4866e0c0",
  1409 => x"02a866c4",
  1410 => x"c487c8c0",
  1411 => x"78c048a6",
  1412 => x"c487c5c0",
  1413 => x"78c148a6",
  1414 => x"c01e66c4",
  1415 => x"49751ee0",
  1416 => x"87ced8ff",
  1417 => x"4c7086c8",
  1418 => x"06acb7c0",
  1419 => x"7487d4c1",
  1420 => x"49e0c085",
  1421 => x"4b758974",
  1422 => x"4ac0ddc1",
  1423 => x"e6e9fe71",
  1424 => x"c085c287",
  1425 => x"c14866e4",
  1426 => x"a6e8c080",
  1427 => x"66ecc058",
  1428 => x"7081c149",
  1429 => x"c8c002a9",
  1430 => x"48a6c487",
  1431 => x"c5c078c0",
  1432 => x"48a6c487",
  1433 => x"66c478c1",
  1434 => x"49a4c21e",
  1435 => x"7148e0c0",
  1436 => x"1e497088",
  1437 => x"d6ff4975",
  1438 => x"86c887f8",
  1439 => x"01a8b7c0",
  1440 => x"c087c0ff",
  1441 => x"c00266e4",
  1442 => x"496e87d1",
  1443 => x"e4c081c9",
  1444 => x"486e5166",
  1445 => x"78ffc6c1",
  1446 => x"6e87ccc0",
  1447 => x"c281c949",
  1448 => x"c1486e51",
  1449 => x"c878eec8",
  1450 => x"66cc4866",
  1451 => x"cbc004a8",
  1452 => x"4866c887",
  1453 => x"a6cc80c1",
  1454 => x"87e9c058",
  1455 => x"c14866cc",
  1456 => x"58a6d088",
  1457 => x"ff87dec0",
  1458 => x"7087d3d5",
  1459 => x"87d5c04c",
  1460 => x"05acc6c1",
  1461 => x"d087c8c0",
  1462 => x"80c14866",
  1463 => x"ff58a6d4",
  1464 => x"7087fbd4",
  1465 => x"4866d44c",
  1466 => x"a6d880c1",
  1467 => x"029c7458",
  1468 => x"c887cbc0",
  1469 => x"c8c14866",
  1470 => x"f204a866",
  1471 => x"d4ff87e8",
  1472 => x"66c887d3",
  1473 => x"03a8c748",
  1474 => x"c287e5c0",
  1475 => x"c048fcef",
  1476 => x"4966c878",
  1477 => x"c0c191cb",
  1478 => x"a1c48166",
  1479 => x"c04a6a4a",
  1480 => x"66c87952",
  1481 => x"cc80c148",
  1482 => x"a8c758a6",
  1483 => x"87dbff04",
  1484 => x"ff8ed0ff",
  1485 => x"4c87e5de",
  1486 => x"2064616f",
  1487 => x"00202e2a",
  1488 => x"1e00203a",
  1489 => x"4b711e73",
  1490 => x"87c6029b",
  1491 => x"48f8efc2",
  1492 => x"1ec778c0",
  1493 => x"bff8efc2",
  1494 => x"e1c11e49",
  1495 => x"efc21ed0",
  1496 => x"ed49bfe0",
  1497 => x"86cc87e8",
  1498 => x"bfe0efc2",
  1499 => x"87e7e849",
  1500 => x"c8029b73",
  1501 => x"d0e1c187",
  1502 => x"c6e3c049",
  1503 => x"dfddff87",
  1504 => x"1e731e87",
  1505 => x"e0c14bc0",
  1506 => x"50c048fc",
  1507 => x"bff3e2c1",
  1508 => x"d9d8ff49",
  1509 => x"05987087",
  1510 => x"dec187c4",
  1511 => x"48734be4",
  1512 => x"87fcdcff",
  1513 => x"204d4f52",
  1514 => x"64616f6c",
  1515 => x"20676e69",
  1516 => x"6c696166",
  1517 => x"1e006465",
  1518 => x"c187dfc7",
  1519 => x"87c3fe49",
  1520 => x"87c9edfe",
  1521 => x"cd029870",
  1522 => x"e2f4fe87",
  1523 => x"02987087",
  1524 => x"4ac187c4",
  1525 => x"4ac087c2",
  1526 => x"ce059a72",
  1527 => x"c11ec087",
  1528 => x"c049c7e0",
  1529 => x"c487d3ee",
  1530 => x"c087fe86",
  1531 => x"d2e0c11e",
  1532 => x"c5eec049",
  1533 => x"fe1ec087",
  1534 => x"497087c7",
  1535 => x"87faedc0",
  1536 => x"f887d6c3",
  1537 => x"534f268e",
  1538 => x"61662044",
  1539 => x"64656c69",
  1540 => x"6f42002e",
  1541 => x"6e69746f",
  1542 => x"2e2e2e67",
  1543 => x"e5c01e00",
  1544 => x"87fa87df",
  1545 => x"c21e4f26",
  1546 => x"c048f8ef",
  1547 => x"e0efc278",
  1548 => x"fe78c048",
  1549 => x"87e587c1",
  1550 => x"4f2648c0",
  1551 => x"00010000",
  1552 => x"20800000",
  1553 => x"74697845",
  1554 => x"42208000",
  1555 => x"006b6361",
  1556 => x"00000f32",
  1557 => x"00002c0c",
  1558 => x"32000000",
  1559 => x"2a00000f",
  1560 => x"0000002c",
  1561 => x"0f320000",
  1562 => x"2c480000",
  1563 => x"00000000",
  1564 => x"000f3200",
  1565 => x"002c6600",
  1566 => x"00000000",
  1567 => x"00000f32",
  1568 => x"00002c84",
  1569 => x"32000000",
  1570 => x"a200000f",
  1571 => x"0000002c",
  1572 => x"0f320000",
  1573 => x"2cc00000",
  1574 => x"00000000",
  1575 => x"00116f00",
  1576 => x"00000000",
  1577 => x"00000000",
  1578 => x"0000123f",
  1579 => x"00000000",
  1580 => x"b7000000",
  1581 => x"50000018",
  1582 => x"30325445",
  1583 => x"52203130",
  1584 => x"1e004d4f",
  1585 => x"c048f0fe",
  1586 => x"7909cd78",
  1587 => x"1e4f2609",
  1588 => x"bff0fe1e",
  1589 => x"2626487e",
  1590 => x"f0fe1e4f",
  1591 => x"2678c148",
  1592 => x"f0fe1e4f",
  1593 => x"2678c048",
  1594 => x"4a711e4f",
  1595 => x"265252c0",
  1596 => x"5b5e0e4f",
  1597 => x"f40e5d5c",
  1598 => x"974d7186",
  1599 => x"a5c17e6d",
  1600 => x"486c974c",
  1601 => x"6e58a6c8",
  1602 => x"a866c448",
  1603 => x"ff87c505",
  1604 => x"87e6c048",
  1605 => x"c287caff",
  1606 => x"6c9749a5",
  1607 => x"4ba3714b",
  1608 => x"974b6b97",
  1609 => x"486e7e6c",
  1610 => x"a6c880c1",
  1611 => x"cc98c758",
  1612 => x"977058a6",
  1613 => x"87e1fe7c",
  1614 => x"8ef44873",
  1615 => x"4c264d26",
  1616 => x"4f264b26",
  1617 => x"5c5b5e0e",
  1618 => x"7186f40e",
  1619 => x"4a66d84c",
  1620 => x"c29affc3",
  1621 => x"6c974ba4",
  1622 => x"49a17349",
  1623 => x"6c975172",
  1624 => x"c1486e7e",
  1625 => x"58a6c880",
  1626 => x"a6cc98c7",
  1627 => x"f4547058",
  1628 => x"87caff8e",
  1629 => x"e8fd1e1e",
  1630 => x"4abfe087",
  1631 => x"c0e0c049",
  1632 => x"87cb0299",
  1633 => x"f3c21e72",
  1634 => x"f7fe49de",
  1635 => x"fc86c487",
  1636 => x"7e7087fd",
  1637 => x"2687c2fd",
  1638 => x"c21e4f26",
  1639 => x"fd49def3",
  1640 => x"e5c187c7",
  1641 => x"dafc49f4",
  1642 => x"87eec387",
  1643 => x"5e0e4f26",
  1644 => x"0e5d5c5b",
  1645 => x"f3c24d71",
  1646 => x"f4fc49de",
  1647 => x"c04b7087",
  1648 => x"c304abb7",
  1649 => x"f0c387c2",
  1650 => x"87c905ab",
  1651 => x"48d2eac1",
  1652 => x"e3c278c1",
  1653 => x"abe0c387",
  1654 => x"c187c905",
  1655 => x"c148d6ea",
  1656 => x"87d4c278",
  1657 => x"bfd6eac1",
  1658 => x"c287c602",
  1659 => x"c24ca3c0",
  1660 => x"c14c7387",
  1661 => x"02bfd2ea",
  1662 => x"7487e0c0",
  1663 => x"29b7c449",
  1664 => x"e9ebc191",
  1665 => x"cf4a7481",
  1666 => x"c192c29a",
  1667 => x"70307248",
  1668 => x"72baff4a",
  1669 => x"70986948",
  1670 => x"7487db79",
  1671 => x"29b7c449",
  1672 => x"e9ebc191",
  1673 => x"cf4a7481",
  1674 => x"c392c29a",
  1675 => x"70307248",
  1676 => x"b069484a",
  1677 => x"9d757970",
  1678 => x"87f0c005",
  1679 => x"c848d0ff",
  1680 => x"d4ff78e1",
  1681 => x"c178c548",
  1682 => x"02bfd6ea",
  1683 => x"e0c387c3",
  1684 => x"d2eac178",
  1685 => x"87c602bf",
  1686 => x"c348d4ff",
  1687 => x"d4ff78f0",
  1688 => x"ff787348",
  1689 => x"e1c848d0",
  1690 => x"78e0c078",
  1691 => x"48d6eac1",
  1692 => x"eac178c0",
  1693 => x"78c048d2",
  1694 => x"49def3c2",
  1695 => x"7087f2f9",
  1696 => x"abb7c04b",
  1697 => x"87fefc03",
  1698 => x"4d2648c0",
  1699 => x"4b264c26",
  1700 => x"00004f26",
  1701 => x"00000000",
  1702 => x"c01e0000",
  1703 => x"c449724a",
  1704 => x"e9ebc191",
  1705 => x"c179c081",
  1706 => x"aab7d082",
  1707 => x"2687ee04",
  1708 => x"5b5e0e4f",
  1709 => x"710e5d5c",
  1710 => x"87e5f84d",
  1711 => x"b7c44a75",
  1712 => x"ebc1922a",
  1713 => x"4c7582e9",
  1714 => x"94c29ccf",
  1715 => x"744b496a",
  1716 => x"c29bc32b",
  1717 => x"70307448",
  1718 => x"74bcff4c",
  1719 => x"70987148",
  1720 => x"87f5f77a",
  1721 => x"e1fe4873",
  1722 => x"00000087",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000000",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"d0ff1e00",
  1739 => x"78e1c848",
  1740 => x"d4ff4871",
  1741 => x"66c47808",
  1742 => x"08d4ff48",
  1743 => x"1e4f2678",
  1744 => x"66c44a71",
  1745 => x"49721e49",
  1746 => x"ff87deff",
  1747 => x"e0c048d0",
  1748 => x"4f262678",
  1749 => x"711e731e",
  1750 => x"4966c84b",
  1751 => x"c14a731e",
  1752 => x"ff49a2e0",
  1753 => x"c42687d9",
  1754 => x"264d2687",
  1755 => x"264b264c",
  1756 => x"d4ff1e4f",
  1757 => x"7affc34a",
  1758 => x"c048d0ff",
  1759 => x"7ade78e1",
  1760 => x"bfe8f3c2",
  1761 => x"c848497a",
  1762 => x"717a7028",
  1763 => x"7028d048",
  1764 => x"d848717a",
  1765 => x"ff7a7028",
  1766 => x"e0c048d0",
  1767 => x"1e4f2678",
  1768 => x"c848d0ff",
  1769 => x"487178c9",
  1770 => x"7808d4ff",
  1771 => x"711e4f26",
  1772 => x"87eb494a",
  1773 => x"c848d0ff",
  1774 => x"1e4f2678",
  1775 => x"4b711e73",
  1776 => x"bff8f3c2",
  1777 => x"c287c302",
  1778 => x"d0ff87eb",
  1779 => x"78c9c848",
  1780 => x"e0c04973",
  1781 => x"48d4ffb1",
  1782 => x"f3c27871",
  1783 => x"78c048ec",
  1784 => x"c50266c8",
  1785 => x"49ffc387",
  1786 => x"49c087c2",
  1787 => x"59f4f3c2",
  1788 => x"c60266cc",
  1789 => x"d5d5c587",
  1790 => x"cf87c44a",
  1791 => x"c24affff",
  1792 => x"c25af8f3",
  1793 => x"c148f8f3",
  1794 => x"2687c478",
  1795 => x"264c264d",
  1796 => x"0e4f264b",
  1797 => x"5d5c5b5e",
  1798 => x"c24a710e",
  1799 => x"4cbff4f3",
  1800 => x"cb029a72",
  1801 => x"91c84987",
  1802 => x"4bf1eec1",
  1803 => x"87c48371",
  1804 => x"4bf1f2c1",
  1805 => x"49134dc0",
  1806 => x"f3c29974",
  1807 => x"ffb9bff0",
  1808 => x"787148d4",
  1809 => x"852cb7c1",
  1810 => x"04adb7c8",
  1811 => x"f3c287e8",
  1812 => x"c848bfec",
  1813 => x"f0f3c280",
  1814 => x"87effe58",
  1815 => x"711e731e",
  1816 => x"9a4a134b",
  1817 => x"7287cb02",
  1818 => x"87e7fe49",
  1819 => x"059a4a13",
  1820 => x"dafe87f5",
  1821 => x"f3c21e87",
  1822 => x"c249bfec",
  1823 => x"c148ecf3",
  1824 => x"c0c478a1",
  1825 => x"db03a9b7",
  1826 => x"48d4ff87",
  1827 => x"bff0f3c2",
  1828 => x"ecf3c278",
  1829 => x"f3c249bf",
  1830 => x"a1c148ec",
  1831 => x"b7c0c478",
  1832 => x"87e504a9",
  1833 => x"c848d0ff",
  1834 => x"f8f3c278",
  1835 => x"2678c048",
  1836 => x"0000004f",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00005f5f",
  1840 => x"03030000",
  1841 => x"00030300",
  1842 => x"7f7f1400",
  1843 => x"147f7f14",
  1844 => x"2e240000",
  1845 => x"123a6b6b",
  1846 => x"366a4c00",
  1847 => x"32566c18",
  1848 => x"4f7e3000",
  1849 => x"683a7759",
  1850 => x"04000040",
  1851 => x"00000307",
  1852 => x"1c000000",
  1853 => x"0041633e",
  1854 => x"41000000",
  1855 => x"001c3e63",
  1856 => x"3e2a0800",
  1857 => x"2a3e1c1c",
  1858 => x"08080008",
  1859 => x"08083e3e",
  1860 => x"80000000",
  1861 => x"000060e0",
  1862 => x"08080000",
  1863 => x"08080808",
  1864 => x"00000000",
  1865 => x"00006060",
  1866 => x"30604000",
  1867 => x"03060c18",
  1868 => x"7f3e0001",
  1869 => x"3e7f4d59",
  1870 => x"06040000",
  1871 => x"00007f7f",
  1872 => x"63420000",
  1873 => x"464f5971",
  1874 => x"63220000",
  1875 => x"367f4949",
  1876 => x"161c1800",
  1877 => x"107f7f13",
  1878 => x"67270000",
  1879 => x"397d4545",
  1880 => x"7e3c0000",
  1881 => x"3079494b",
  1882 => x"01010000",
  1883 => x"070f7971",
  1884 => x"7f360000",
  1885 => x"367f4949",
  1886 => x"4f060000",
  1887 => x"1e3f6949",
  1888 => x"00000000",
  1889 => x"00006666",
  1890 => x"80000000",
  1891 => x"000066e6",
  1892 => x"08080000",
  1893 => x"22221414",
  1894 => x"14140000",
  1895 => x"14141414",
  1896 => x"22220000",
  1897 => x"08081414",
  1898 => x"03020000",
  1899 => x"060f5951",
  1900 => x"417f3e00",
  1901 => x"1e1f555d",
  1902 => x"7f7e0000",
  1903 => x"7e7f0909",
  1904 => x"7f7f0000",
  1905 => x"367f4949",
  1906 => x"3e1c0000",
  1907 => x"41414163",
  1908 => x"7f7f0000",
  1909 => x"1c3e6341",
  1910 => x"7f7f0000",
  1911 => x"41414949",
  1912 => x"7f7f0000",
  1913 => x"01010909",
  1914 => x"7f3e0000",
  1915 => x"7a7b4941",
  1916 => x"7f7f0000",
  1917 => x"7f7f0808",
  1918 => x"41000000",
  1919 => x"00417f7f",
  1920 => x"60200000",
  1921 => x"3f7f4040",
  1922 => x"087f7f00",
  1923 => x"4163361c",
  1924 => x"7f7f0000",
  1925 => x"40404040",
  1926 => x"067f7f00",
  1927 => x"7f7f060c",
  1928 => x"067f7f00",
  1929 => x"7f7f180c",
  1930 => x"7f3e0000",
  1931 => x"3e7f4141",
  1932 => x"7f7f0000",
  1933 => x"060f0909",
  1934 => x"417f3e00",
  1935 => x"407e7f61",
  1936 => x"7f7f0000",
  1937 => x"667f1909",
  1938 => x"6f260000",
  1939 => x"327b594d",
  1940 => x"01010000",
  1941 => x"01017f7f",
  1942 => x"7f3f0000",
  1943 => x"3f7f4040",
  1944 => x"3f0f0000",
  1945 => x"0f3f7070",
  1946 => x"307f7f00",
  1947 => x"7f7f3018",
  1948 => x"36634100",
  1949 => x"63361c1c",
  1950 => x"06030141",
  1951 => x"03067c7c",
  1952 => x"59716101",
  1953 => x"4143474d",
  1954 => x"7f000000",
  1955 => x"0041417f",
  1956 => x"06030100",
  1957 => x"6030180c",
  1958 => x"41000040",
  1959 => x"007f7f41",
  1960 => x"060c0800",
  1961 => x"080c0603",
  1962 => x"80808000",
  1963 => x"80808080",
  1964 => x"00000000",
  1965 => x"00040703",
  1966 => x"74200000",
  1967 => x"787c5454",
  1968 => x"7f7f0000",
  1969 => x"387c4444",
  1970 => x"7c380000",
  1971 => x"00444444",
  1972 => x"7c380000",
  1973 => x"7f7f4444",
  1974 => x"7c380000",
  1975 => x"185c5454",
  1976 => x"7e040000",
  1977 => x"0005057f",
  1978 => x"bc180000",
  1979 => x"7cfca4a4",
  1980 => x"7f7f0000",
  1981 => x"787c0404",
  1982 => x"00000000",
  1983 => x"00407d3d",
  1984 => x"80800000",
  1985 => x"007dfd80",
  1986 => x"7f7f0000",
  1987 => x"446c3810",
  1988 => x"00000000",
  1989 => x"00407f3f",
  1990 => x"0c7c7c00",
  1991 => x"787c0c18",
  1992 => x"7c7c0000",
  1993 => x"787c0404",
  1994 => x"7c380000",
  1995 => x"387c4444",
  1996 => x"fcfc0000",
  1997 => x"183c2424",
  1998 => x"3c180000",
  1999 => x"fcfc2424",
  2000 => x"7c7c0000",
  2001 => x"080c0404",
  2002 => x"5c480000",
  2003 => x"20745454",
  2004 => x"3f040000",
  2005 => x"0044447f",
  2006 => x"7c3c0000",
  2007 => x"7c7c4040",
  2008 => x"3c1c0000",
  2009 => x"1c3c6060",
  2010 => x"607c3c00",
  2011 => x"3c7c6030",
  2012 => x"386c4400",
  2013 => x"446c3810",
  2014 => x"bc1c0000",
  2015 => x"1c3c60e0",
  2016 => x"64440000",
  2017 => x"444c5c74",
  2018 => x"08080000",
  2019 => x"4141773e",
  2020 => x"00000000",
  2021 => x"00007f7f",
  2022 => x"41410000",
  2023 => x"08083e77",
  2024 => x"01010200",
  2025 => x"01020203",
  2026 => x"7f7f7f00",
  2027 => x"7f7f7f7f",
  2028 => x"1c080800",
  2029 => x"7f3e3e1c",
  2030 => x"3e7f7f7f",
  2031 => x"081c1c3e",
  2032 => x"18100008",
  2033 => x"10187c7c",
  2034 => x"30100000",
  2035 => x"10307c7c",
  2036 => x"60301000",
  2037 => x"061e7860",
  2038 => x"3c664200",
  2039 => x"42663c18",
  2040 => x"6a387800",
  2041 => x"386cc6c2",
  2042 => x"00006000",
  2043 => x"60000060",
  2044 => x"5b5e0e00",
  2045 => x"1e0e5d5c",
  2046 => x"f4c24c71",
  2047 => x"c04dbfc9",
  2048 => x"741ec04b",
  2049 => x"87c702ab",
  2050 => x"c048a6c4",
  2051 => x"c487c578",
  2052 => x"78c148a6",
  2053 => x"731e66c4",
  2054 => x"87dfee49",
  2055 => x"e0c086c8",
  2056 => x"87efef49",
  2057 => x"6a4aa5c4",
  2058 => x"87f0f049",
  2059 => x"cb87c6f1",
  2060 => x"c883c185",
  2061 => x"ff04abb7",
  2062 => x"262687c7",
  2063 => x"264c264d",
  2064 => x"1e4f264b",
  2065 => x"f4c24a71",
  2066 => x"f4c25acd",
  2067 => x"78c748cd",
  2068 => x"87ddfe49",
  2069 => x"731e4f26",
  2070 => x"c04a711e",
  2071 => x"d303aab7",
  2072 => x"d3cfc287",
  2073 => x"87c405bf",
  2074 => x"87c24bc1",
  2075 => x"cfc24bc0",
  2076 => x"87c45bd7",
  2077 => x"5ad7cfc2",
  2078 => x"bfd3cfc2",
  2079 => x"c19ac14a",
  2080 => x"ec49a2c0",
  2081 => x"48fc87e8",
  2082 => x"bfd3cfc2",
  2083 => x"87effe78",
  2084 => x"c44a711e",
  2085 => x"49721e66",
  2086 => x"2687f9ea",
  2087 => x"711e4f26",
  2088 => x"48d4ff4a",
  2089 => x"ff78ffc3",
  2090 => x"e1c048d0",
  2091 => x"48d4ff78",
  2092 => x"497278c1",
  2093 => x"787131c4",
  2094 => x"c048d0ff",
  2095 => x"4f2678e0",
  2096 => x"d3cfc21e",
  2097 => x"cbda49bf",
  2098 => x"c1f4c287",
  2099 => x"78bfe848",
  2100 => x"48fdf3c2",
  2101 => x"c278bfec",
  2102 => x"4abfc1f4",
  2103 => x"99ffc349",
  2104 => x"722ab7c8",
  2105 => x"c2b07148",
  2106 => x"2658c9f4",
  2107 => x"5b5e0e4f",
  2108 => x"710e5d5c",
  2109 => x"87c8ff4b",
  2110 => x"48fcf3c2",
  2111 => x"497350c0",
  2112 => x"7087eee6",
  2113 => x"9cc24c49",
  2114 => x"cb49eecb",
  2115 => x"497087cd",
  2116 => x"fcf3c24d",
  2117 => x"c105bf97",
  2118 => x"66d087e2",
  2119 => x"c5f4c249",
  2120 => x"d60599bf",
  2121 => x"4966d487",
  2122 => x"bffdf3c2",
  2123 => x"87cb0599",
  2124 => x"fce54973",
  2125 => x"02987087",
  2126 => x"c187c1c1",
  2127 => x"87c0fe4c",
  2128 => x"e2ca4975",
  2129 => x"02987087",
  2130 => x"f3c287c6",
  2131 => x"50c148fc",
  2132 => x"97fcf3c2",
  2133 => x"e3c005bf",
  2134 => x"c5f4c287",
  2135 => x"66d049bf",
  2136 => x"d6ff0599",
  2137 => x"fdf3c287",
  2138 => x"66d449bf",
  2139 => x"caff0599",
  2140 => x"e4497387",
  2141 => x"987087fb",
  2142 => x"87fffe05",
  2143 => x"fafa4874",
  2144 => x"5b5e0e87",
  2145 => x"f80e5d5c",
  2146 => x"4c4dc086",
  2147 => x"c47ebfec",
  2148 => x"f4c248a6",
  2149 => x"c178bfc9",
  2150 => x"c71ec01e",
  2151 => x"87cdfd49",
  2152 => x"987086c8",
  2153 => x"ff87cd02",
  2154 => x"87eafa49",
  2155 => x"e349dac1",
  2156 => x"4dc187ff",
  2157 => x"97fcf3c2",
  2158 => x"87cf02bf",
  2159 => x"bfcbcfc2",
  2160 => x"c2b9c149",
  2161 => x"7159cfcf",
  2162 => x"c287d3fb",
  2163 => x"4bbfc1f4",
  2164 => x"bfd3cfc2",
  2165 => x"87e9c005",
  2166 => x"e349fdc3",
  2167 => x"fac387d3",
  2168 => x"87cde349",
  2169 => x"ffc34973",
  2170 => x"c01e7199",
  2171 => x"87e0fa49",
  2172 => x"b7c84973",
  2173 => x"c11e7129",
  2174 => x"87d4fa49",
  2175 => x"f4c586c8",
  2176 => x"c5f4c287",
  2177 => x"029b4bbf",
  2178 => x"cfc287dd",
  2179 => x"c749bfcf",
  2180 => x"987087d5",
  2181 => x"c087c405",
  2182 => x"c287d24b",
  2183 => x"fac649e0",
  2184 => x"d3cfc287",
  2185 => x"c287c658",
  2186 => x"c048cfcf",
  2187 => x"c2497378",
  2188 => x"87cd0599",
  2189 => x"e149ebc3",
  2190 => x"497087f7",
  2191 => x"c20299c2",
  2192 => x"734cfb87",
  2193 => x"0599c149",
  2194 => x"f4c387cd",
  2195 => x"87e1e149",
  2196 => x"99c24970",
  2197 => x"fa87c202",
  2198 => x"c849734c",
  2199 => x"87cd0599",
  2200 => x"e149f5c3",
  2201 => x"497087cb",
  2202 => x"d50299c2",
  2203 => x"cdf4c287",
  2204 => x"87ca02bf",
  2205 => x"c288c148",
  2206 => x"c058d1f4",
  2207 => x"4cff87c2",
  2208 => x"49734dc1",
  2209 => x"cd0599c4",
  2210 => x"49f2c387",
  2211 => x"7087e2e0",
  2212 => x"0299c249",
  2213 => x"f4c287dc",
  2214 => x"487ebfcd",
  2215 => x"03a8b7c7",
  2216 => x"6e87cbc0",
  2217 => x"c280c148",
  2218 => x"c058d1f4",
  2219 => x"4cfe87c2",
  2220 => x"fdc34dc1",
  2221 => x"f8dfff49",
  2222 => x"c2497087",
  2223 => x"87d50299",
  2224 => x"bfcdf4c2",
  2225 => x"87c9c002",
  2226 => x"48cdf4c2",
  2227 => x"c2c078c0",
  2228 => x"c14cfd87",
  2229 => x"49fac34d",
  2230 => x"87d5dfff",
  2231 => x"99c24970",
  2232 => x"87d9c002",
  2233 => x"bfcdf4c2",
  2234 => x"a8b7c748",
  2235 => x"87c9c003",
  2236 => x"48cdf4c2",
  2237 => x"c2c078c7",
  2238 => x"c14cfc87",
  2239 => x"acb7c04d",
  2240 => x"87d3c003",
  2241 => x"c14866c4",
  2242 => x"7e7080d8",
  2243 => x"c002bf6e",
  2244 => x"744b87c5",
  2245 => x"c00f7349",
  2246 => x"1ef0c31e",
  2247 => x"f749dac1",
  2248 => x"86c887cb",
  2249 => x"c0029870",
  2250 => x"f4c287d8",
  2251 => x"6e7ebfcd",
  2252 => x"c491cb49",
  2253 => x"82714a66",
  2254 => x"c5c0026a",
  2255 => x"496e4b87",
  2256 => x"9d750f73",
  2257 => x"87c8c002",
  2258 => x"bfcdf4c2",
  2259 => x"87e1f249",
  2260 => x"bfd7cfc2",
  2261 => x"87ddc002",
  2262 => x"87cbc249",
  2263 => x"c0029870",
  2264 => x"f4c287d3",
  2265 => x"f249bfcd",
  2266 => x"49c087c7",
  2267 => x"c287e7f3",
  2268 => x"c048d7cf",
  2269 => x"f38ef878",
  2270 => x"5e0e87c1",
  2271 => x"0e5d5c5b",
  2272 => x"c24c711e",
  2273 => x"49bfc9f4",
  2274 => x"4da1cdc1",
  2275 => x"6981d1c1",
  2276 => x"029c747e",
  2277 => x"a5c487cf",
  2278 => x"c27b744b",
  2279 => x"49bfc9f4",
  2280 => x"6e87e0f2",
  2281 => x"059c747b",
  2282 => x"4bc087c4",
  2283 => x"4bc187c2",
  2284 => x"e1f24973",
  2285 => x"0266d487",
  2286 => x"de4987c7",
  2287 => x"c24a7087",
  2288 => x"c24ac087",
  2289 => x"265adbcf",
  2290 => x"0087f0f1",
  2291 => x"00000000",
  2292 => x"00000000",
  2293 => x"00000000",
  2294 => x"1e000000",
  2295 => x"c8ff4a71",
  2296 => x"a17249bf",
  2297 => x"1e4f2648",
  2298 => x"89bfc8ff",
  2299 => x"c0c0c0fe",
  2300 => x"01a9c0c0",
  2301 => x"4ac087c4",
  2302 => x"4ac187c2",
  2303 => x"4f264872",
  2304 => x"dcd3ff1e",
  2305 => x"4966c487",
  2306 => x"0299c0c2",
  2307 => x"e0c387cd",
  2308 => x"def3c21e",
  2309 => x"ebd4ff49",
  2310 => x"c486c487",
  2311 => x"c0c44966",
  2312 => x"87cd0299",
  2313 => x"c21ef0c3",
  2314 => x"ff49def3",
  2315 => x"c487d5d4",
  2316 => x"4966c486",
  2317 => x"7199ffc1",
  2318 => x"def3c21e",
  2319 => x"c3d4ff49",
  2320 => x"d4d2ff87",
  2321 => x"4f262687",
  2322 => x"5c5b5e0e",
  2323 => x"dcff0e5d",
  2324 => x"c27ec086",
  2325 => x"49bfd5f4",
  2326 => x"1e7181c2",
  2327 => x"4ac61e72",
  2328 => x"87c7f2fd",
  2329 => x"4a264871",
  2330 => x"a6c84926",
  2331 => x"d5f4c258",
  2332 => x"81c449bf",
  2333 => x"1e721e71",
  2334 => x"f1fd4ac6",
  2335 => x"487187ed",
  2336 => x"49264a26",
  2337 => x"c258a6cc",
  2338 => x"49bfeedc",
  2339 => x"7087d8fd",
  2340 => x"ceca0298",
  2341 => x"49e0c087",
  2342 => x"7087c0fd",
  2343 => x"f2dcc249",
  2344 => x"744cc059",
  2345 => x"fe91c449",
  2346 => x"4a6981d0",
  2347 => x"f4c24974",
  2348 => x"c481bfd5",
  2349 => x"e5f4c291",
  2350 => x"9a797281",
  2351 => x"7287d202",
  2352 => x"7189c149",
  2353 => x"c1486e9a",
  2354 => x"727e7080",
  2355 => x"eeff059a",
  2356 => x"c284c187",
  2357 => x"ff04acb7",
  2358 => x"486e87c9",
  2359 => x"a8b7fcc0",
  2360 => x"87ffc804",
  2361 => x"4a744cc0",
  2362 => x"c48266c4",
  2363 => x"e5f4c292",
  2364 => x"c8497482",
  2365 => x"91c48166",
  2366 => x"81e5f4c2",
  2367 => x"49694a6a",
  2368 => x"4b74b972",
  2369 => x"bfd5f4c2",
  2370 => x"c293c483",
  2371 => x"6b83e5f4",
  2372 => x"714872ba",
  2373 => x"58a6d098",
  2374 => x"f4c24974",
  2375 => x"c481bfd5",
  2376 => x"e5f4c291",
  2377 => x"d07e6981",
  2378 => x"78c048a6",
  2379 => x"df4966cc",
  2380 => x"c0c70229",
  2381 => x"c04a7487",
  2382 => x"66d092e0",
  2383 => x"48ffc082",
  2384 => x"4a708872",
  2385 => x"c048a6d4",
  2386 => x"c080c478",
  2387 => x"df496e78",
  2388 => x"a6e0c029",
  2389 => x"d1f4c259",
  2390 => x"7278c148",
  2391 => x"b731c349",
  2392 => x"c0b1722a",
  2393 => x"91c499ff",
  2394 => x"4dc5dec2",
  2395 => x"4b6d8571",
  2396 => x"c0c0c449",
  2397 => x"f3c00299",
  2398 => x"0266dc87",
  2399 => x"80c887c8",
  2400 => x"c57840c0",
  2401 => x"f4c287ef",
  2402 => x"78c148d9",
  2403 => x"bfddf4c2",
  2404 => x"87e1c505",
  2405 => x"f81ed8c1",
  2406 => x"e3f949a0",
  2407 => x"1ed8c587",
  2408 => x"49d1f4c2",
  2409 => x"c887d9f9",
  2410 => x"87c9c586",
  2411 => x"d80266dc",
  2412 => x"c2497387",
  2413 => x"0299c0c0",
  2414 => x"d087c3c0",
  2415 => x"486d2bb7",
  2416 => x"98fffffd",
  2417 => x"fac07d70",
  2418 => x"d9f4c287",
  2419 => x"f2c002bf",
  2420 => x"d0487387",
  2421 => x"e4c028b7",
  2422 => x"987058a6",
  2423 => x"87e3c002",
  2424 => x"bfe1f4c2",
  2425 => x"c0e0c049",
  2426 => x"cac00299",
  2427 => x"c0497087",
  2428 => x"0299c0e0",
  2429 => x"6d87ccc0",
  2430 => x"c0c0c248",
  2431 => x"c07d70b0",
  2432 => x"734b66e0",
  2433 => x"c0c0c849",
  2434 => x"c7c20299",
  2435 => x"e1f4c287",
  2436 => x"c0cc4abf",
  2437 => x"cfc0029a",
  2438 => x"8ac0c487",
  2439 => x"87d8c002",
  2440 => x"f9c0028a",
  2441 => x"87ddc187",
  2442 => x"ffc34973",
  2443 => x"c291c299",
  2444 => x"1181f9dd",
  2445 => x"87dcc14b",
  2446 => x"ffc34973",
  2447 => x"c291c299",
  2448 => x"c181f9dd",
  2449 => x"dc4b1181",
  2450 => x"c8c00266",
  2451 => x"48a6d887",
  2452 => x"ffc078d2",
  2453 => x"48a6d487",
  2454 => x"c078d2c4",
  2455 => x"497387f6",
  2456 => x"c299ffc3",
  2457 => x"f9ddc291",
  2458 => x"1181c181",
  2459 => x"0266dc4b",
  2460 => x"d887c9c0",
  2461 => x"d9c148a6",
  2462 => x"87d8c078",
  2463 => x"c548a6d4",
  2464 => x"cfc078d9",
  2465 => x"c3497387",
  2466 => x"91c299ff",
  2467 => x"81f9ddc2",
  2468 => x"4b1181c1",
  2469 => x"c00266dc",
  2470 => x"497387dc",
  2471 => x"fcc7b9ff",
  2472 => x"487199c0",
  2473 => x"bfe1f4c2",
  2474 => x"e5f4c298",
  2475 => x"9bffc358",
  2476 => x"c0b3c0c4",
  2477 => x"497387d4",
  2478 => x"99c0fcc7",
  2479 => x"f4c24871",
  2480 => x"c2b0bfe1",
  2481 => x"c358e5f4",
  2482 => x"66d49bff",
  2483 => x"87cac002",
  2484 => x"d1f4c21e",
  2485 => x"87e8f449",
  2486 => x"1e7386c4",
  2487 => x"49d1f4c2",
  2488 => x"c487ddf4",
  2489 => x"0266d886",
  2490 => x"1e87cac0",
  2491 => x"49d1f4c2",
  2492 => x"c487cdf4",
  2493 => x"4866cc86",
  2494 => x"a6d030c1",
  2495 => x"c1486e58",
  2496 => x"d07e7030",
  2497 => x"80c14866",
  2498 => x"c058a6d4",
  2499 => x"04a8b7e0",
  2500 => x"c187d9f8",
  2501 => x"acb7c284",
  2502 => x"87caf704",
  2503 => x"48d5f4c2",
  2504 => x"ff7866c4",
  2505 => x"4d268edc",
  2506 => x"4b264c26",
  2507 => x"00004f26",
  2508 => x"c01e0000",
  2509 => x"c449724a",
  2510 => x"e5f4c291",
  2511 => x"c179ff81",
  2512 => x"aab7c682",
  2513 => x"c287ee04",
  2514 => x"c048d5f4",
  2515 => x"80c87840",
  2516 => x"4f2678c0",
  2517 => x"711e731e",
  2518 => x"f5ddc24b",
  2519 => x"87c905bf",
  2520 => x"48f5ddc2",
  2521 => x"c9ff78c1",
  2522 => x"87dcf387",
  2523 => x"c8ff4973",
  2524 => x"f5fe87fc",
  2525 => x"00000087",
  2526 => x"f2ebf400",
  2527 => x"040605f5",
  2528 => x"830b030c",
  2529 => x"fc00660a",
  2530 => x"da005a00",
  2531 => x"94800000",
  2532 => x"78800508",
  2533 => x"01800200",
  2534 => x"09800300",
  2535 => x"00800400",
  2536 => x"91800100",
  2537 => x"04002608",
  2538 => x"00001d00",
  2539 => x"00001c00",
  2540 => x"0c002500",
  2541 => x"00001a00",
  2542 => x"00001b00",
  2543 => x"00002400",
  2544 => x"00011200",
  2545 => x"03002e00",
  2546 => x"00002d00",
  2547 => x"00002300",
  2548 => x"0b003600",
  2549 => x"00002100",
  2550 => x"00002b00",
  2551 => x"00002c00",
  2552 => x"00002200",
  2553 => x"6c003d00",
  2554 => x"00003500",
  2555 => x"00003400",
  2556 => x"75003e00",
  2557 => x"00003200",
  2558 => x"00003300",
  2559 => x"6b003c00",
  2560 => x"00002a00",
  2561 => x"01004600",
  2562 => x"73004300",
  2563 => x"69003b00",
  2564 => x"09004500",
  2565 => x"70003a00",
  2566 => x"72004200",
  2567 => x"74004400",
  2568 => x"00003100",
  2569 => x"00005500",
  2570 => x"7c004d00",
  2571 => x"7a004b00",
  2572 => x"00007b00",
  2573 => x"71004900",
  2574 => x"84004c00",
  2575 => x"77005400",
  2576 => x"00004100",
  2577 => x"00006100",
  2578 => x"7c005b00",
  2579 => x"00005200",
  2580 => x"0000f100",
  2581 => x"00025900",
  2582 => x"5d000e00",
  2583 => x"00005d00",
  2584 => x"79004a00",
  2585 => x"05001600",
  2586 => x"07007600",
  2587 => x"0d000d00",
  2588 => x"06001e00",
  2589 => x"00002900",
  2590 => x"00041400",
  2591 => x"00001500",
  2592 => x"00400000",
  2593 => x"00400000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
