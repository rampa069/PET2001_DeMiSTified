library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"4c711e0e",
     1 => x"bfd1f4c2",
     2 => x"c04bc04d",
     3 => x"02ab741e",
     4 => x"a6c487c7",
     5 => x"c578c048",
     6 => x"48a6c487",
     7 => x"66c478c1",
     8 => x"ee49731e",
     9 => x"86c887df",
    10 => x"ef49e0c0",
    11 => x"a5c487ef",
    12 => x"f0496a4a",
    13 => x"c6f187f0",
    14 => x"c185cb87",
    15 => x"abb7c883",
    16 => x"87c7ff04",
    17 => x"264d2626",
    18 => x"264b264c",
    19 => x"4a711e4f",
    20 => x"5ad5f4c2",
    21 => x"48d5f4c2",
    22 => x"fe4978c7",
    23 => x"4f2687dd",
    24 => x"711e731e",
    25 => x"aab7c04a",
    26 => x"c287d303",
    27 => x"05bfdecf",
    28 => x"4bc187c4",
    29 => x"4bc087c2",
    30 => x"5be2cfc2",
    31 => x"cfc287c4",
    32 => x"cfc25ae2",
    33 => x"c14abfde",
    34 => x"a2c0c19a",
    35 => x"87e8ec49",
    36 => x"cfc248fc",
    37 => x"fe78bfde",
    38 => x"711e87ef",
    39 => x"1e66c44a",
    40 => x"f9e94972",
    41 => x"4f262687",
    42 => x"ff4a711e",
    43 => x"ffc348d4",
    44 => x"48d0ff78",
    45 => x"ff78e1c0",
    46 => x"78c148d4",
    47 => x"31c44972",
    48 => x"d0ff7871",
    49 => x"78e0c048",
    50 => x"c21e4f26",
    51 => x"49bfdecf",
    52 => x"c287ccda",
    53 => x"e848c9f4",
    54 => x"f4c278bf",
    55 => x"bfec48c5",
    56 => x"c9f4c278",
    57 => x"c3494abf",
    58 => x"b7c899ff",
    59 => x"7148722a",
    60 => x"d1f4c2b0",
    61 => x"0e4f2658",
    62 => x"5d5c5b5e",
    63 => x"ff4b710e",
    64 => x"f4c287c8",
    65 => x"50c048c4",
    66 => x"eee54973",
    67 => x"4c497087",
    68 => x"eecb9cc2",
    69 => x"87cecb49",
    70 => x"c24d4970",
    71 => x"bf97c4f4",
    72 => x"87e2c105",
    73 => x"c24966d0",
    74 => x"99bfcdf4",
    75 => x"d487d605",
    76 => x"f4c24966",
    77 => x"0599bfc5",
    78 => x"497387cb",
    79 => x"7087fce4",
    80 => x"c1c10298",
    81 => x"fe4cc187",
    82 => x"497587c0",
    83 => x"7087e3ca",
    84 => x"87c60298",
    85 => x"48c4f4c2",
    86 => x"f4c250c1",
    87 => x"05bf97c4",
    88 => x"c287e3c0",
    89 => x"49bfcdf4",
    90 => x"059966d0",
    91 => x"c287d6ff",
    92 => x"49bfc5f4",
    93 => x"059966d4",
    94 => x"7387caff",
    95 => x"87fbe349",
    96 => x"fe059870",
    97 => x"487487ff",
    98 => x"0e87fafa",
    99 => x"5d5c5b5e",
   100 => x"c086f80e",
   101 => x"bfec4c4d",
   102 => x"48a6c47e",
   103 => x"bfd1f4c2",
   104 => x"c01ec178",
   105 => x"fd49c71e",
   106 => x"86c887cd",
   107 => x"cd029870",
   108 => x"fa49ff87",
   109 => x"dac187ea",
   110 => x"87ffe249",
   111 => x"f4c24dc1",
   112 => x"02bf97c4",
   113 => x"cfc287cf",
   114 => x"c149bfd6",
   115 => x"dacfc2b9",
   116 => x"d3fb7159",
   117 => x"c9f4c287",
   118 => x"cfc24bbf",
   119 => x"c005bfde",
   120 => x"fdc387e9",
   121 => x"87d3e249",
   122 => x"e249fac3",
   123 => x"497387cd",
   124 => x"7199ffc3",
   125 => x"fa49c01e",
   126 => x"497387e0",
   127 => x"7129b7c8",
   128 => x"fa49c11e",
   129 => x"86c887d4",
   130 => x"c287f5c5",
   131 => x"4bbfcdf4",
   132 => x"87dd029b",
   133 => x"bfdacfc2",
   134 => x"87d6c749",
   135 => x"c4059870",
   136 => x"d24bc087",
   137 => x"49e0c287",
   138 => x"c287fbc6",
   139 => x"c658decf",
   140 => x"dacfc287",
   141 => x"7378c048",
   142 => x"0599c249",
   143 => x"ebc387cd",
   144 => x"87f7e049",
   145 => x"99c24970",
   146 => x"fb87c202",
   147 => x"c149734c",
   148 => x"87cd0599",
   149 => x"e049f4c3",
   150 => x"497087e1",
   151 => x"c20299c2",
   152 => x"734cfa87",
   153 => x"0599c849",
   154 => x"f5c387cd",
   155 => x"87cbe049",
   156 => x"99c24970",
   157 => x"c287d502",
   158 => x"02bfd5f4",
   159 => x"c14887ca",
   160 => x"d9f4c288",
   161 => x"87c2c058",
   162 => x"4dc14cff",
   163 => x"99c44973",
   164 => x"c387ce05",
   165 => x"dfff49f2",
   166 => x"497087e1",
   167 => x"dc0299c2",
   168 => x"d5f4c287",
   169 => x"c7487ebf",
   170 => x"c003a8b7",
   171 => x"486e87cb",
   172 => x"f4c280c1",
   173 => x"c2c058d9",
   174 => x"c14cfe87",
   175 => x"49fdc34d",
   176 => x"87f7deff",
   177 => x"99c24970",
   178 => x"c287d502",
   179 => x"02bfd5f4",
   180 => x"c287c9c0",
   181 => x"c048d5f4",
   182 => x"87c2c078",
   183 => x"4dc14cfd",
   184 => x"ff49fac3",
   185 => x"7087d4de",
   186 => x"0299c249",
   187 => x"c287d9c0",
   188 => x"48bfd5f4",
   189 => x"03a8b7c7",
   190 => x"c287c9c0",
   191 => x"c748d5f4",
   192 => x"87c2c078",
   193 => x"4dc14cfc",
   194 => x"03acb7c0",
   195 => x"c487d3c0",
   196 => x"d8c14866",
   197 => x"6e7e7080",
   198 => x"c5c002bf",
   199 => x"49744b87",
   200 => x"1ec00f73",
   201 => x"c11ef0c3",
   202 => x"caf749da",
   203 => x"7086c887",
   204 => x"d8c00298",
   205 => x"d5f4c287",
   206 => x"496e7ebf",
   207 => x"66c491cb",
   208 => x"6a82714a",
   209 => x"87c5c002",
   210 => x"73496e4b",
   211 => x"029d750f",
   212 => x"c287c8c0",
   213 => x"49bfd5f4",
   214 => x"c287e0f2",
   215 => x"02bfe2cf",
   216 => x"4987ddc0",
   217 => x"7087cbc2",
   218 => x"d3c00298",
   219 => x"d5f4c287",
   220 => x"c6f249bf",
   221 => x"f349c087",
   222 => x"cfc287e6",
   223 => x"78c048e2",
   224 => x"c0f38ef8",
   225 => x"5b5e0e87",
   226 => x"1e0e5d5c",
   227 => x"f4c24c71",
   228 => x"c149bfd1",
   229 => x"c14da1cd",
   230 => x"7e6981d1",
   231 => x"cf029c74",
   232 => x"4ba5c487",
   233 => x"f4c27b74",
   234 => x"f249bfd1",
   235 => x"7b6e87df",
   236 => x"c4059c74",
   237 => x"c24bc087",
   238 => x"734bc187",
   239 => x"87e0f249",
   240 => x"c70266d4",
   241 => x"87de4987",
   242 => x"87c24a70",
   243 => x"cfc24ac0",
   244 => x"f1265ae6",
   245 => x"000087ef",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"00000000",
   249 => x"711e0000",
   250 => x"bfc8ff4a",
   251 => x"48a17249",
   252 => x"ff1e4f26",
   253 => x"fe89bfc8",
   254 => x"c0c0c0c0",
   255 => x"c401a9c0",
   256 => x"c24ac087",
   257 => x"724ac187",
   258 => x"1e4f2648",
   259 => x"87dbd2ff",
   260 => x"c24966c4",
   261 => x"cd0299c0",
   262 => x"1ee0c387",
   263 => x"49e6f3c2",
   264 => x"87ead3ff",
   265 => x"66c486c4",
   266 => x"99c0c449",
   267 => x"c387cd02",
   268 => x"f3c21ef0",
   269 => x"d3ff49e6",
   270 => x"86c487d4",
   271 => x"c14966c4",
   272 => x"1e7199ff",
   273 => x"49e6f3c2",
   274 => x"87c2d3ff",
   275 => x"87d3d1ff",
   276 => x"0e4f2626",
   277 => x"5d5c5b5e",
   278 => x"86dcff0e",
   279 => x"f4c27ec0",
   280 => x"c249bfdd",
   281 => x"721e7181",
   282 => x"fd4ac61e",
   283 => x"7187fcf1",
   284 => x"264a2648",
   285 => x"58a6c849",
   286 => x"bfddf4c2",
   287 => x"7181c449",
   288 => x"c61e721e",
   289 => x"e2f1fd4a",
   290 => x"26487187",
   291 => x"cc49264a",
   292 => x"dcc258a6",
   293 => x"fd49bff9",
   294 => x"987087d8",
   295 => x"87ceca02",
   296 => x"fd49e0c0",
   297 => x"497087c0",
   298 => x"59fddcc2",
   299 => x"49744cc0",
   300 => x"d0fe91c4",
   301 => x"744a6981",
   302 => x"ddf4c249",
   303 => x"91c481bf",
   304 => x"81edf4c2",
   305 => x"029a7972",
   306 => x"497287d2",
   307 => x"9a7189c1",
   308 => x"80c1486e",
   309 => x"9a727e70",
   310 => x"87eeff05",
   311 => x"b7c284c1",
   312 => x"c9ff04ac",
   313 => x"c0486e87",
   314 => x"04a8b7fc",
   315 => x"c087ffc8",
   316 => x"c44a744c",
   317 => x"92c48266",
   318 => x"82edf4c2",
   319 => x"66c84974",
   320 => x"c291c481",
   321 => x"6a81edf4",
   322 => x"7249694a",
   323 => x"c24b74b9",
   324 => x"83bfddf4",
   325 => x"f4c293c4",
   326 => x"ba6b83ed",
   327 => x"98714872",
   328 => x"7458a6d0",
   329 => x"ddf4c249",
   330 => x"91c481bf",
   331 => x"81edf4c2",
   332 => x"a6d07e69",
   333 => x"cc78c048",
   334 => x"29df4966",
   335 => x"87c0c702",
   336 => x"e0c04a74",
   337 => x"8266d092",
   338 => x"7248ffc0",
   339 => x"d44a7088",
   340 => x"78c048a6",
   341 => x"78c080c4",
   342 => x"29df496e",
   343 => x"59a6e0c0",
   344 => x"48d9f4c2",
   345 => x"497278c1",
   346 => x"2ab731c3",
   347 => x"ffc0b172",
   348 => x"c291c499",
   349 => x"714dd0de",
   350 => x"494b6d85",
   351 => x"99c0c0c4",
   352 => x"87f3c002",
   353 => x"c80266dc",
   354 => x"c080c887",
   355 => x"efc57840",
   356 => x"e1f4c287",
   357 => x"c278c148",
   358 => x"05bfe5f4",
   359 => x"c187e1c5",
   360 => x"a0f81ed8",
   361 => x"87e3f949",
   362 => x"c21ed8c5",
   363 => x"f949d9f4",
   364 => x"86c887d9",
   365 => x"dc87c9c5",
   366 => x"87d80266",
   367 => x"c0c24973",
   368 => x"c00299c0",
   369 => x"b7d087c3",
   370 => x"fd486d2b",
   371 => x"7098ffff",
   372 => x"87fac07d",
   373 => x"bfe1f4c2",
   374 => x"87f2c002",
   375 => x"b7d04873",
   376 => x"a6e4c028",
   377 => x"02987058",
   378 => x"c287e3c0",
   379 => x"49bfe9f4",
   380 => x"99c0e0c0",
   381 => x"87cac002",
   382 => x"e0c04970",
   383 => x"c00299c0",
   384 => x"486d87cc",
   385 => x"b0c0c0c2",
   386 => x"e0c07d70",
   387 => x"49734b66",
   388 => x"99c0c0c8",
   389 => x"87c7c202",
   390 => x"bfe9f4c2",
   391 => x"9ac0cc4a",
   392 => x"87cfc002",
   393 => x"028ac0c4",
   394 => x"8a87d8c0",
   395 => x"87f9c002",
   396 => x"7387ddc1",
   397 => x"99ffc349",
   398 => x"dec291c2",
   399 => x"4b1181c4",
   400 => x"7387dcc1",
   401 => x"99ffc349",
   402 => x"dec291c2",
   403 => x"81c181c4",
   404 => x"66dc4b11",
   405 => x"87c8c002",
   406 => x"d248a6d8",
   407 => x"87ffc078",
   408 => x"c448a6d4",
   409 => x"f6c078d2",
   410 => x"c3497387",
   411 => x"91c299ff",
   412 => x"81c4dec2",
   413 => x"4b1181c1",
   414 => x"c00266dc",
   415 => x"a6d887c9",
   416 => x"78d9c148",
   417 => x"d487d8c0",
   418 => x"d9c548a6",
   419 => x"87cfc078",
   420 => x"ffc34973",
   421 => x"c291c299",
   422 => x"c181c4de",
   423 => x"dc4b1181",
   424 => x"dcc00266",
   425 => x"ff497387",
   426 => x"c0fcc7b9",
   427 => x"c2487199",
   428 => x"98bfe9f4",
   429 => x"58edf4c2",
   430 => x"c49bffc3",
   431 => x"d4c0b3c0",
   432 => x"c7497387",
   433 => x"7199c0fc",
   434 => x"e9f4c248",
   435 => x"f4c2b0bf",
   436 => x"ffc358ed",
   437 => x"0266d49b",
   438 => x"1e87cac0",
   439 => x"49d9f4c2",
   440 => x"c487e8f4",
   441 => x"c21e7386",
   442 => x"f449d9f4",
   443 => x"86c487dd",
   444 => x"c00266d8",
   445 => x"c21e87ca",
   446 => x"f449d9f4",
   447 => x"86c487cd",
   448 => x"c14866cc",
   449 => x"58a6d030",
   450 => x"30c1486e",
   451 => x"66d07e70",
   452 => x"d480c148",
   453 => x"e0c058a6",
   454 => x"f804a8b7",
   455 => x"84c187d9",
   456 => x"04acb7c2",
   457 => x"c287caf7",
   458 => x"c448ddf4",
   459 => x"dcff7866",
   460 => x"264d268e",
   461 => x"264b264c",
   462 => x"0000004f",
   463 => x"4ac01e00",
   464 => x"91c44972",
   465 => x"81edf4c2",
   466 => x"82c179ff",
   467 => x"04aab7c6",
   468 => x"f4c287ee",
   469 => x"40c048dd",
   470 => x"c080c878",
   471 => x"1e4f2678",
   472 => x"4b711e73",
   473 => x"bfc0dec2",
   474 => x"c287c905",
   475 => x"c148c0de",
   476 => x"87c9ff78",
   477 => x"7387dcf3",
   478 => x"fbc7ff49",
   479 => x"87f5fe87",
   480 => x"00000000",
   481 => x"f5f2ebf4",
   482 => x"0c040605",
   483 => x"0a830b03",
   484 => x"00fc0066",
   485 => x"00da005a",
   486 => x"08948000",
   487 => x"00788005",
   488 => x"00018002",
   489 => x"00098003",
   490 => x"00008004",
   491 => x"08918001",
   492 => x"00040026",
   493 => x"0000001d",
   494 => x"0000001c",
   495 => x"000c0025",
   496 => x"0000001a",
   497 => x"0000001b",
   498 => x"00000024",
   499 => x"00000112",
   500 => x"0003002e",
   501 => x"0000002d",
   502 => x"00000023",
   503 => x"000b0036",
   504 => x"00000021",
   505 => x"0000002b",
   506 => x"0000002c",
   507 => x"00000022",
   508 => x"006c003d",
   509 => x"00000035",
   510 => x"00000034",
   511 => x"0075003e",
   512 => x"00000032",
   513 => x"00000033",
   514 => x"006b003c",
   515 => x"0000002a",
   516 => x"00010046",
   517 => x"00730043",
   518 => x"0069003b",
   519 => x"00090045",
   520 => x"0070003a",
   521 => x"00720042",
   522 => x"00740044",
   523 => x"00000031",
   524 => x"00000055",
   525 => x"007c004d",
   526 => x"007a004b",
   527 => x"0000007b",
   528 => x"00710049",
   529 => x"0084004c",
   530 => x"00770054",
   531 => x"00000041",
   532 => x"00000061",
   533 => x"007c005b",
   534 => x"00000052",
   535 => x"000000f1",
   536 => x"00000259",
   537 => x"005d000e",
   538 => x"0000005d",
   539 => x"0079004a",
   540 => x"00050016",
   541 => x"00070076",
   542 => x"000d000d",
   543 => x"0006001e",
   544 => x"00000029",
   545 => x"00000414",
   546 => x"00000015",
   547 => x"00004000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
