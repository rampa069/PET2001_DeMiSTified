library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e0f5c287",
    12 => x"86c0c84e",
    13 => x"49e0f5c2",
    14 => x"48d0e2c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e5de",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"9a721e73",
    47 => x"87e7c002",
    48 => x"4bc148c0",
    49 => x"d106a972",
    50 => x"06827287",
    51 => x"837387c9",
    52 => x"f401a972",
    53 => x"c187c387",
    54 => x"a9723ab2",
    55 => x"80738903",
    56 => x"2b2ac107",
    57 => x"2687f305",
    58 => x"1e4f264b",
    59 => x"4dc41e75",
    60 => x"04a1b771",
    61 => x"81c1b9ff",
    62 => x"7207bdc3",
    63 => x"ff04a2b7",
    64 => x"c182c1ba",
    65 => x"eefe07bd",
    66 => x"042dc187",
    67 => x"80c1b8ff",
    68 => x"ff042d07",
    69 => x"0781c1b9",
    70 => x"4f264d26",
    71 => x"c44a711e",
    72 => x"c1484966",
    73 => x"58a6c888",
    74 => x"d6029971",
    75 => x"48d4ff87",
    76 => x"6878ffc3",
    77 => x"4966c452",
    78 => x"c888c148",
    79 => x"997158a6",
    80 => x"2687ea05",
    81 => x"1e731e4f",
    82 => x"c34bd4ff",
    83 => x"4a6b7bff",
    84 => x"6b7bffc3",
    85 => x"7232c849",
    86 => x"7bffc3b1",
    87 => x"31c84a6b",
    88 => x"ffc3b271",
    89 => x"c8496b7b",
    90 => x"71b17232",
    91 => x"2687c448",
    92 => x"264c264d",
    93 => x"0e4f264b",
    94 => x"5d5c5b5e",
    95 => x"ff4a710e",
    96 => x"49724cd4",
    97 => x"7199ffc3",
    98 => x"d0e2c27c",
    99 => x"87c805bf",
   100 => x"c94866d0",
   101 => x"58a6d430",
   102 => x"d84966d0",
   103 => x"99ffc329",
   104 => x"66d07c71",
   105 => x"c329d049",
   106 => x"7c7199ff",
   107 => x"c84966d0",
   108 => x"99ffc329",
   109 => x"66d07c71",
   110 => x"99ffc349",
   111 => x"49727c71",
   112 => x"ffc329d0",
   113 => x"6c7c7199",
   114 => x"fff0c94b",
   115 => x"abffc34d",
   116 => x"c387d005",
   117 => x"4b6c7cff",
   118 => x"c6028dc1",
   119 => x"abffc387",
   120 => x"7387f002",
   121 => x"87c7fe48",
   122 => x"ff49c01e",
   123 => x"ffc348d4",
   124 => x"c381c178",
   125 => x"04a9b7c8",
   126 => x"4f2687f1",
   127 => x"e71e731e",
   128 => x"dff8c487",
   129 => x"c01ec04b",
   130 => x"f7c1f0ff",
   131 => x"87e7fd49",
   132 => x"a8c186c4",
   133 => x"87eac005",
   134 => x"c348d4ff",
   135 => x"c0c178ff",
   136 => x"c0c0c0c0",
   137 => x"f0e1c01e",
   138 => x"fd49e9c1",
   139 => x"86c487c9",
   140 => x"ca059870",
   141 => x"48d4ff87",
   142 => x"c178ffc3",
   143 => x"fe87cb48",
   144 => x"8bc187e6",
   145 => x"87fdfe05",
   146 => x"e6fc48c0",
   147 => x"1e731e87",
   148 => x"c348d4ff",
   149 => x"4bd378ff",
   150 => x"ffc01ec0",
   151 => x"49c1c1f0",
   152 => x"c487d4fc",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187f1fd",
   158 => x"dbff058b",
   159 => x"fb48c087",
   160 => x"5e0e87f1",
   161 => x"ff0e5c5b",
   162 => x"dbfd4cd4",
   163 => x"1eeac687",
   164 => x"c1f0e1c0",
   165 => x"defb49c8",
   166 => x"c186c487",
   167 => x"87c802a8",
   168 => x"c087eafe",
   169 => x"87e2c148",
   170 => x"7087dafa",
   171 => x"ffffcf49",
   172 => x"a9eac699",
   173 => x"fe87c802",
   174 => x"48c087d3",
   175 => x"c387cbc1",
   176 => x"f1c07cff",
   177 => x"87f4fc4b",
   178 => x"c0029870",
   179 => x"1ec087eb",
   180 => x"c1f0ffc0",
   181 => x"defa49fa",
   182 => x"7086c487",
   183 => x"87d90598",
   184 => x"6c7cffc3",
   185 => x"7cffc349",
   186 => x"c17c7c7c",
   187 => x"c40299c0",
   188 => x"d548c187",
   189 => x"d148c087",
   190 => x"05abc287",
   191 => x"48c087c4",
   192 => x"8bc187c8",
   193 => x"87fdfe05",
   194 => x"e4f948c0",
   195 => x"1e731e87",
   196 => x"48d0e2c2",
   197 => x"4bc778c1",
   198 => x"c248d0ff",
   199 => x"87c8fb78",
   200 => x"c348d0ff",
   201 => x"c01ec078",
   202 => x"c0c1d0e5",
   203 => x"87c7f949",
   204 => x"a8c186c4",
   205 => x"4b87c105",
   206 => x"c505abc2",
   207 => x"c048c087",
   208 => x"8bc187f9",
   209 => x"87d0ff05",
   210 => x"c287f7fc",
   211 => x"7058d4e2",
   212 => x"87cd0598",
   213 => x"ffc01ec1",
   214 => x"49d0c1f0",
   215 => x"c487d8f8",
   216 => x"48d4ff86",
   217 => x"c278ffc3",
   218 => x"e2c287fc",
   219 => x"d0ff58d8",
   220 => x"ff78c248",
   221 => x"ffc348d4",
   222 => x"f748c178",
   223 => x"5e0e87f5",
   224 => x"0e5d5c5b",
   225 => x"4cc04b71",
   226 => x"dfcdeec5",
   227 => x"48d4ff4a",
   228 => x"6878ffc3",
   229 => x"a9fec349",
   230 => x"87fdc005",
   231 => x"9b734d70",
   232 => x"d087cc02",
   233 => x"49731e66",
   234 => x"c487f1f5",
   235 => x"ff87d686",
   236 => x"d1c448d0",
   237 => x"7dffc378",
   238 => x"c14866d0",
   239 => x"58a6d488",
   240 => x"f0059870",
   241 => x"48d4ff87",
   242 => x"7878ffc3",
   243 => x"c5059b73",
   244 => x"48d0ff87",
   245 => x"4ac178d0",
   246 => x"058ac14c",
   247 => x"7487eefe",
   248 => x"87cbf648",
   249 => x"711e731e",
   250 => x"ff4bc04a",
   251 => x"ffc348d4",
   252 => x"48d0ff78",
   253 => x"ff78c3c4",
   254 => x"ffc348d4",
   255 => x"c01e7278",
   256 => x"d1c1f0ff",
   257 => x"87eff549",
   258 => x"987086c4",
   259 => x"c887d205",
   260 => x"66cc1ec0",
   261 => x"87e6fd49",
   262 => x"4b7086c4",
   263 => x"c248d0ff",
   264 => x"f5487378",
   265 => x"5e0e87cd",
   266 => x"0e5d5c5b",
   267 => x"ffc01ec0",
   268 => x"49c9c1f0",
   269 => x"d287c0f5",
   270 => x"d8e2c21e",
   271 => x"87fefc49",
   272 => x"4cc086c8",
   273 => x"b7d284c1",
   274 => x"87f804ac",
   275 => x"97d8e2c2",
   276 => x"c0c349bf",
   277 => x"a9c0c199",
   278 => x"87e7c005",
   279 => x"97dfe2c2",
   280 => x"31d049bf",
   281 => x"97e0e2c2",
   282 => x"32c84abf",
   283 => x"e2c2b172",
   284 => x"4abf97e1",
   285 => x"cf4c71b1",
   286 => x"9cffffff",
   287 => x"34ca84c1",
   288 => x"c287e7c1",
   289 => x"bf97e1e2",
   290 => x"c631c149",
   291 => x"e2e2c299",
   292 => x"c74abf97",
   293 => x"b1722ab7",
   294 => x"97dde2c2",
   295 => x"cf4d4abf",
   296 => x"dee2c29d",
   297 => x"c34abf97",
   298 => x"c232ca9a",
   299 => x"bf97dfe2",
   300 => x"7333c24b",
   301 => x"e0e2c2b2",
   302 => x"c34bbf97",
   303 => x"b7c69bc0",
   304 => x"c2b2732b",
   305 => x"7148c181",
   306 => x"c1497030",
   307 => x"70307548",
   308 => x"c14c724d",
   309 => x"c8947184",
   310 => x"06adb7c0",
   311 => x"34c187cc",
   312 => x"c0c82db7",
   313 => x"ff01adb7",
   314 => x"487487f4",
   315 => x"0e87c0f2",
   316 => x"5d5c5b5e",
   317 => x"c286f80e",
   318 => x"c048feea",
   319 => x"f6e2c278",
   320 => x"fb49c01e",
   321 => x"86c487de",
   322 => x"c5059870",
   323 => x"c948c087",
   324 => x"4dc087ce",
   325 => x"efc07ec1",
   326 => x"c249bfd8",
   327 => x"714aece3",
   328 => x"c4ed4bc8",
   329 => x"05987087",
   330 => x"7ec087c2",
   331 => x"bfd4efc0",
   332 => x"c8e4c249",
   333 => x"4bc8714a",
   334 => x"7087eeec",
   335 => x"87c20598",
   336 => x"026e7ec0",
   337 => x"c287fdc0",
   338 => x"4dbffce9",
   339 => x"9ff4eac2",
   340 => x"c5487ebf",
   341 => x"05a8ead6",
   342 => x"e9c287c7",
   343 => x"ce4dbffc",
   344 => x"ca486e87",
   345 => x"02a8d5e9",
   346 => x"48c087c5",
   347 => x"c287f1c7",
   348 => x"751ef6e2",
   349 => x"87ecf949",
   350 => x"987086c4",
   351 => x"c087c505",
   352 => x"87dcc748",
   353 => x"bfd4efc0",
   354 => x"c8e4c249",
   355 => x"4bc8714a",
   356 => x"7087d6eb",
   357 => x"87c80598",
   358 => x"48feeac2",
   359 => x"87da78c1",
   360 => x"bfd8efc0",
   361 => x"ece3c249",
   362 => x"4bc8714a",
   363 => x"7087faea",
   364 => x"c5c00298",
   365 => x"c648c087",
   366 => x"eac287e6",
   367 => x"49bf97f4",
   368 => x"05a9d5c1",
   369 => x"c287cdc0",
   370 => x"bf97f5ea",
   371 => x"a9eac249",
   372 => x"87c5c002",
   373 => x"c7c648c0",
   374 => x"f6e2c287",
   375 => x"487ebf97",
   376 => x"02a8e9c3",
   377 => x"6e87cec0",
   378 => x"a8ebc348",
   379 => x"87c5c002",
   380 => x"ebc548c0",
   381 => x"c1e3c287",
   382 => x"9949bf97",
   383 => x"87ccc005",
   384 => x"97c2e3c2",
   385 => x"a9c249bf",
   386 => x"87c5c002",
   387 => x"cfc548c0",
   388 => x"c3e3c287",
   389 => x"c248bf97",
   390 => x"7058faea",
   391 => x"88c1484c",
   392 => x"58feeac2",
   393 => x"97c4e3c2",
   394 => x"817549bf",
   395 => x"97c5e3c2",
   396 => x"32c84abf",
   397 => x"c27ea172",
   398 => x"6e48cbef",
   399 => x"c6e3c278",
   400 => x"c848bf97",
   401 => x"eac258a6",
   402 => x"c202bffe",
   403 => x"efc087d4",
   404 => x"c249bfd4",
   405 => x"714ac8e4",
   406 => x"cce84bc8",
   407 => x"02987087",
   408 => x"c087c5c0",
   409 => x"87f8c348",
   410 => x"bff6eac2",
   411 => x"dfefc24c",
   412 => x"dbe3c25c",
   413 => x"c849bf97",
   414 => x"dae3c231",
   415 => x"a14abf97",
   416 => x"dce3c249",
   417 => x"d04abf97",
   418 => x"49a17232",
   419 => x"97dde3c2",
   420 => x"32d84abf",
   421 => x"c449a172",
   422 => x"efc29166",
   423 => x"c281bfcb",
   424 => x"c259d3ef",
   425 => x"bf97e3e3",
   426 => x"c232c84a",
   427 => x"bf97e2e3",
   428 => x"c24aa24b",
   429 => x"bf97e4e3",
   430 => x"7333d04b",
   431 => x"e3c24aa2",
   432 => x"4bbf97e5",
   433 => x"33d89bcf",
   434 => x"c24aa273",
   435 => x"c25ad7ef",
   436 => x"4abfd3ef",
   437 => x"92748ac2",
   438 => x"48d7efc2",
   439 => x"c178a172",
   440 => x"e3c287ca",
   441 => x"49bf97c8",
   442 => x"e3c231c8",
   443 => x"4abf97c7",
   444 => x"ebc249a1",
   445 => x"ebc259c6",
   446 => x"c549bfc2",
   447 => x"81ffc731",
   448 => x"efc229c9",
   449 => x"e3c259df",
   450 => x"4abf97cd",
   451 => x"e3c232c8",
   452 => x"4bbf97cc",
   453 => x"66c44aa2",
   454 => x"c2826e92",
   455 => x"c25adbef",
   456 => x"c048d3ef",
   457 => x"cfefc278",
   458 => x"78a17248",
   459 => x"48dfefc2",
   460 => x"bfd3efc2",
   461 => x"e3efc278",
   462 => x"d7efc248",
   463 => x"eac278bf",
   464 => x"c002bffe",
   465 => x"487487c9",
   466 => x"7e7030c4",
   467 => x"c287c9c0",
   468 => x"48bfdbef",
   469 => x"7e7030c4",
   470 => x"48c2ebc2",
   471 => x"48c1786e",
   472 => x"4d268ef8",
   473 => x"4b264c26",
   474 => x"5e0e4f26",
   475 => x"0e5d5c5b",
   476 => x"eac24a71",
   477 => x"cb02bffe",
   478 => x"c74b7287",
   479 => x"c14c722b",
   480 => x"87c99cff",
   481 => x"2bc84b72",
   482 => x"ffc34c72",
   483 => x"cbefc29c",
   484 => x"efc083bf",
   485 => x"02abbfd0",
   486 => x"efc087d9",
   487 => x"e2c25bd4",
   488 => x"49731ef6",
   489 => x"c487fdf0",
   490 => x"05987086",
   491 => x"48c087c5",
   492 => x"c287e6c0",
   493 => x"02bffeea",
   494 => x"497487d2",
   495 => x"e2c291c4",
   496 => x"4d6981f6",
   497 => x"ffffffcf",
   498 => x"87cb9dff",
   499 => x"91c24974",
   500 => x"81f6e2c2",
   501 => x"754d699f",
   502 => x"87c6fe48",
   503 => x"5c5b5e0e",
   504 => x"86f80e5d",
   505 => x"059c4c71",
   506 => x"48c087c5",
   507 => x"c887c2c3",
   508 => x"486e7ea4",
   509 => x"66d878c0",
   510 => x"d887c702",
   511 => x"05bf9766",
   512 => x"48c087c5",
   513 => x"c087eac2",
   514 => x"4949c11e",
   515 => x"c487e6c7",
   516 => x"9d4d7086",
   517 => x"87c2c102",
   518 => x"4ac6ebc2",
   519 => x"e04966d8",
   520 => x"987087ec",
   521 => x"87f2c002",
   522 => x"66d84a75",
   523 => x"e14bcb49",
   524 => x"987087d1",
   525 => x"87e2c002",
   526 => x"9d751ec0",
   527 => x"c887c702",
   528 => x"78c048a6",
   529 => x"a6c887c5",
   530 => x"c878c148",
   531 => x"e4c64966",
   532 => x"7086c487",
   533 => x"fe059d4d",
   534 => x"9d7587fe",
   535 => x"87cfc102",
   536 => x"6e49a5dc",
   537 => x"da786948",
   538 => x"a6c449a5",
   539 => x"78a4c448",
   540 => x"c448699f",
   541 => x"c2780866",
   542 => x"02bffeea",
   543 => x"a5d487d2",
   544 => x"49699f49",
   545 => x"99ffffc0",
   546 => x"30d04871",
   547 => x"87c27e70",
   548 => x"496e7ec0",
   549 => x"bf66c448",
   550 => x"0866c480",
   551 => x"cc7cc078",
   552 => x"66c449a4",
   553 => x"a4d079bf",
   554 => x"c179c049",
   555 => x"c087c248",
   556 => x"fa8ef848",
   557 => x"5e0e87ec",
   558 => x"0e5d5c5b",
   559 => x"029c4c71",
   560 => x"c887cac1",
   561 => x"026949a4",
   562 => x"d087c2c1",
   563 => x"496c4a66",
   564 => x"5aa6d482",
   565 => x"b94d66d0",
   566 => x"bffaeac2",
   567 => x"72baff4a",
   568 => x"02997199",
   569 => x"c487e4c0",
   570 => x"496b4ba4",
   571 => x"7087fbf9",
   572 => x"f6eac27b",
   573 => x"816c49bf",
   574 => x"b9757c71",
   575 => x"bffaeac2",
   576 => x"72baff4a",
   577 => x"05997199",
   578 => x"7587dcff",
   579 => x"87d2f97c",
   580 => x"711e731e",
   581 => x"c7029b4b",
   582 => x"49a3c887",
   583 => x"87c50569",
   584 => x"f7c048c0",
   585 => x"cfefc287",
   586 => x"a3c44abf",
   587 => x"c2496949",
   588 => x"f6eac289",
   589 => x"a27191bf",
   590 => x"faeac24a",
   591 => x"996b49bf",
   592 => x"c04aa271",
   593 => x"c85ad4ef",
   594 => x"49721e66",
   595 => x"c487d5ea",
   596 => x"05987086",
   597 => x"48c087c4",
   598 => x"48c187c2",
   599 => x"1e87c7f8",
   600 => x"4b711e73",
   601 => x"e4c0029b",
   602 => x"e3efc287",
   603 => x"c24a735b",
   604 => x"f6eac28a",
   605 => x"c29249bf",
   606 => x"48bfcfef",
   607 => x"efc28072",
   608 => x"487158e7",
   609 => x"ebc230c4",
   610 => x"edc058c6",
   611 => x"dfefc287",
   612 => x"d3efc248",
   613 => x"efc278bf",
   614 => x"efc248e3",
   615 => x"c278bfd7",
   616 => x"02bffeea",
   617 => x"eac287c9",
   618 => x"c449bff6",
   619 => x"c287c731",
   620 => x"49bfdbef",
   621 => x"ebc231c4",
   622 => x"e9f659c6",
   623 => x"5b5e0e87",
   624 => x"4a710e5c",
   625 => x"9a724bc0",
   626 => x"87e1c002",
   627 => x"9f49a2da",
   628 => x"eac24b69",
   629 => x"cf02bffe",
   630 => x"49a2d487",
   631 => x"4c49699f",
   632 => x"9cffffc0",
   633 => x"87c234d0",
   634 => x"49744cc0",
   635 => x"fd4973b3",
   636 => x"eff587ed",
   637 => x"5b5e0e87",
   638 => x"f40e5d5c",
   639 => x"c04a7186",
   640 => x"029a727e",
   641 => x"e2c287d8",
   642 => x"78c048f2",
   643 => x"48eae2c2",
   644 => x"bfe3efc2",
   645 => x"eee2c278",
   646 => x"dfefc248",
   647 => x"ebc278bf",
   648 => x"50c048d3",
   649 => x"bfc2ebc2",
   650 => x"f2e2c249",
   651 => x"aa714abf",
   652 => x"87c9c403",
   653 => x"99cf4972",
   654 => x"87e9c005",
   655 => x"48d0efc0",
   656 => x"bfeae2c2",
   657 => x"f6e2c278",
   658 => x"eae2c21e",
   659 => x"e2c249bf",
   660 => x"a1c148ea",
   661 => x"cbe67178",
   662 => x"c086c487",
   663 => x"c248ccef",
   664 => x"cc78f6e2",
   665 => x"ccefc087",
   666 => x"e0c048bf",
   667 => x"d0efc080",
   668 => x"f2e2c258",
   669 => x"80c148bf",
   670 => x"58f6e2c2",
   671 => x"000bcc27",
   672 => x"bf97bf00",
   673 => x"c2029d4d",
   674 => x"e5c387e3",
   675 => x"dcc202ad",
   676 => x"ccefc087",
   677 => x"a3cb4bbf",
   678 => x"cf4c1149",
   679 => x"d2c105ac",
   680 => x"df497587",
   681 => x"cd89c199",
   682 => x"c6ebc291",
   683 => x"4aa3c181",
   684 => x"a3c35112",
   685 => x"c551124a",
   686 => x"51124aa3",
   687 => x"124aa3c7",
   688 => x"4aa3c951",
   689 => x"a3ce5112",
   690 => x"d051124a",
   691 => x"51124aa3",
   692 => x"124aa3d2",
   693 => x"4aa3d451",
   694 => x"a3d65112",
   695 => x"d851124a",
   696 => x"51124aa3",
   697 => x"124aa3dc",
   698 => x"4aa3de51",
   699 => x"7ec15112",
   700 => x"7487fac0",
   701 => x"0599c849",
   702 => x"7487ebc0",
   703 => x"0599d049",
   704 => x"66dc87d1",
   705 => x"87cbc002",
   706 => x"66dc4973",
   707 => x"0298700f",
   708 => x"6e87d3c0",
   709 => x"87c6c005",
   710 => x"48c6ebc2",
   711 => x"efc050c0",
   712 => x"c248bfcc",
   713 => x"ebc287e1",
   714 => x"50c048d3",
   715 => x"c2ebc27e",
   716 => x"e2c249bf",
   717 => x"714abff2",
   718 => x"f7fb04aa",
   719 => x"e3efc287",
   720 => x"c8c005bf",
   721 => x"feeac287",
   722 => x"f8c102bf",
   723 => x"eee2c287",
   724 => x"d5f049bf",
   725 => x"c2497087",
   726 => x"c459f2e2",
   727 => x"e2c248a6",
   728 => x"c278bfee",
   729 => x"02bffeea",
   730 => x"c487d8c0",
   731 => x"ffcf4966",
   732 => x"99f8ffff",
   733 => x"c5c002a9",
   734 => x"c04cc087",
   735 => x"4cc187e1",
   736 => x"c487dcc0",
   737 => x"ffcf4966",
   738 => x"02a999f8",
   739 => x"c887c8c0",
   740 => x"78c048a6",
   741 => x"c887c5c0",
   742 => x"78c148a6",
   743 => x"744c66c8",
   744 => x"e0c0059c",
   745 => x"4966c487",
   746 => x"eac289c2",
   747 => x"914abff6",
   748 => x"bfcfefc2",
   749 => x"eae2c24a",
   750 => x"78a17248",
   751 => x"48f2e2c2",
   752 => x"dff978c0",
   753 => x"f448c087",
   754 => x"87d6ee8e",
   755 => x"00000000",
   756 => x"ffffffff",
   757 => x"00000bdc",
   758 => x"00000be5",
   759 => x"33544146",
   760 => x"20202032",
   761 => x"54414600",
   762 => x"20203631",
   763 => x"ff1e0020",
   764 => x"ffc348d4",
   765 => x"26486878",
   766 => x"d4ff1e4f",
   767 => x"78ffc348",
   768 => x"c048d0ff",
   769 => x"d4ff78e1",
   770 => x"c278d448",
   771 => x"ff48e7ef",
   772 => x"2650bfd4",
   773 => x"d0ff1e4f",
   774 => x"78e0c048",
   775 => x"ff1e4f26",
   776 => x"497087cc",
   777 => x"87c60299",
   778 => x"05a9fbc0",
   779 => x"487187f1",
   780 => x"5e0e4f26",
   781 => x"710e5c5b",
   782 => x"fe4cc04b",
   783 => x"497087f0",
   784 => x"f9c00299",
   785 => x"a9ecc087",
   786 => x"87f2c002",
   787 => x"02a9fbc0",
   788 => x"cc87ebc0",
   789 => x"03acb766",
   790 => x"66d087c7",
   791 => x"7187c202",
   792 => x"02997153",
   793 => x"84c187c2",
   794 => x"7087c3fe",
   795 => x"cd029949",
   796 => x"a9ecc087",
   797 => x"c087c702",
   798 => x"ff05a9fb",
   799 => x"66d087d5",
   800 => x"c087c302",
   801 => x"ecc07b97",
   802 => x"87c405a9",
   803 => x"87c54a74",
   804 => x"0ac04a74",
   805 => x"c248728a",
   806 => x"264d2687",
   807 => x"264b264c",
   808 => x"c9fd1e4f",
   809 => x"4a497087",
   810 => x"04aaf0c0",
   811 => x"f9c087c9",
   812 => x"87c301aa",
   813 => x"c18af0c0",
   814 => x"c904aac1",
   815 => x"aadac187",
   816 => x"c087c301",
   817 => x"48728af7",
   818 => x"5e0e4f26",
   819 => x"710e5c5b",
   820 => x"4bd4ff4a",
   821 => x"e7c04972",
   822 => x"9c4c7087",
   823 => x"c187c202",
   824 => x"48d0ff8c",
   825 => x"d5c178c5",
   826 => x"c649747b",
   827 => x"c6e0c131",
   828 => x"484abf97",
   829 => x"7b70b071",
   830 => x"c448d0ff",
   831 => x"87dbfe78",
   832 => x"5c5b5e0e",
   833 => x"86f80e5d",
   834 => x"7ec04c71",
   835 => x"c087eafb",
   836 => x"edf6c04b",
   837 => x"c049bf97",
   838 => x"87cf04a9",
   839 => x"c187fffb",
   840 => x"edf6c083",
   841 => x"ab49bf97",
   842 => x"c087f106",
   843 => x"bf97edf6",
   844 => x"fa87cf02",
   845 => x"497087f8",
   846 => x"87c60299",
   847 => x"05a9ecc0",
   848 => x"4bc087f1",
   849 => x"7087e7fa",
   850 => x"87e2fa4d",
   851 => x"fa58a6c8",
   852 => x"4a7087dc",
   853 => x"a4c883c1",
   854 => x"49699749",
   855 => x"87c702ad",
   856 => x"05adffc0",
   857 => x"c987e7c0",
   858 => x"699749a4",
   859 => x"a966c449",
   860 => x"4887c702",
   861 => x"05a8ffc0",
   862 => x"a4ca87d4",
   863 => x"49699749",
   864 => x"87c602aa",
   865 => x"05aaffc0",
   866 => x"7ec187c4",
   867 => x"ecc087d0",
   868 => x"87c602ad",
   869 => x"05adfbc0",
   870 => x"4bc087c4",
   871 => x"026e7ec1",
   872 => x"f987e1fe",
   873 => x"487387ef",
   874 => x"ecfb8ef8",
   875 => x"5e0e0087",
   876 => x"0e5d5c5b",
   877 => x"4d7186f8",
   878 => x"754bd4ff",
   879 => x"ecefc21e",
   880 => x"87d8e849",
   881 => x"987086c4",
   882 => x"87ccc402",
   883 => x"c148a6c4",
   884 => x"78bfc8e0",
   885 => x"f1fb4975",
   886 => x"48d0ff87",
   887 => x"d6c178c5",
   888 => x"754ac07b",
   889 => x"7b1149a2",
   890 => x"b7cb82c1",
   891 => x"87f304aa",
   892 => x"ffc34acc",
   893 => x"c082c17b",
   894 => x"04aab7e0",
   895 => x"d0ff87f4",
   896 => x"c378c448",
   897 => x"78c57bff",
   898 => x"c17bd3c1",
   899 => x"6678c47b",
   900 => x"a8b7c048",
   901 => x"87f0c206",
   902 => x"bff4efc2",
   903 => x"4866c44c",
   904 => x"a6c88874",
   905 => x"029c7458",
   906 => x"c287f9c1",
   907 => x"c87ef6e2",
   908 => x"c08c4dc0",
   909 => x"c603acb7",
   910 => x"a4c0c887",
   911 => x"c24cc04d",
   912 => x"bf97e7ef",
   913 => x"0299d049",
   914 => x"1ec087d1",
   915 => x"49ecefc2",
   916 => x"c487fdea",
   917 => x"4a497086",
   918 => x"c287eec0",
   919 => x"c21ef6e2",
   920 => x"ea49ecef",
   921 => x"86c487ea",
   922 => x"ff4a4970",
   923 => x"c5c848d0",
   924 => x"7bd4c178",
   925 => x"7bbf976e",
   926 => x"80c1486e",
   927 => x"8dc17e70",
   928 => x"87f0ff05",
   929 => x"c448d0ff",
   930 => x"059a7278",
   931 => x"48c087c5",
   932 => x"c187c7c1",
   933 => x"ecefc21e",
   934 => x"87dae849",
   935 => x"9c7486c4",
   936 => x"87c7fe05",
   937 => x"c04866c4",
   938 => x"d106a8b7",
   939 => x"ecefc287",
   940 => x"d078c048",
   941 => x"f478c080",
   942 => x"f8efc280",
   943 => x"66c478bf",
   944 => x"a8b7c048",
   945 => x"87d0fd01",
   946 => x"c548d0ff",
   947 => x"7bd3c178",
   948 => x"78c47bc0",
   949 => x"87c248c1",
   950 => x"8ef848c0",
   951 => x"4c264d26",
   952 => x"4f264b26",
   953 => x"5c5b5e0e",
   954 => x"711e0e5d",
   955 => x"4d4cc04b",
   956 => x"e8c004ab",
   957 => x"c0f4c087",
   958 => x"029d751e",
   959 => x"4ac087c4",
   960 => x"4ac187c2",
   961 => x"eceb4972",
   962 => x"7086c487",
   963 => x"6e84c17e",
   964 => x"7387c205",
   965 => x"7385c14c",
   966 => x"d8ff06ac",
   967 => x"26486e87",
   968 => x"1e87f9fe",
   969 => x"66c44a71",
   970 => x"7287c505",
   971 => x"87fef949",
   972 => x"5e0e4f26",
   973 => x"0e5d5c5b",
   974 => x"494c711e",
   975 => x"f0c291de",
   976 => x"85714dd4",
   977 => x"c1026d97",
   978 => x"f0c287dd",
   979 => x"744abfc0",
   980 => x"fe497282",
   981 => x"7e7087ce",
   982 => x"c0029848",
   983 => x"f0c287f2",
   984 => x"4a704bc8",
   985 => x"c4ff49cb",
   986 => x"4b7487fd",
   987 => x"e0c193cb",
   988 => x"83c483da",
   989 => x"7bebfec0",
   990 => x"c1c14974",
   991 => x"7b7587fd",
   992 => x"97c7e0c1",
   993 => x"c21e49bf",
   994 => x"fe49c8f0",
   995 => x"86c487d5",
   996 => x"c1c14974",
   997 => x"49c087e5",
   998 => x"87c4c3c1",
   999 => x"48e8efc2",
  1000 => x"49c178c0",
  1001 => x"2687e6dd",
  1002 => x"4c87f1fc",
  1003 => x"6964616f",
  1004 => x"2e2e676e",
  1005 => x"5e0e002e",
  1006 => x"710e5c5b",
  1007 => x"f0c24a4b",
  1008 => x"7282bfc0",
  1009 => x"87dcfc49",
  1010 => x"029c4c70",
  1011 => x"e74987c4",
  1012 => x"f0c287eb",
  1013 => x"78c048c0",
  1014 => x"f0dc49c1",
  1015 => x"87fefb87",
  1016 => x"5c5b5e0e",
  1017 => x"86f40e5d",
  1018 => x"4df6e2c2",
  1019 => x"a6c44cc0",
  1020 => x"c278c048",
  1021 => x"49bfc0f0",
  1022 => x"c106a9c0",
  1023 => x"e2c287c1",
  1024 => x"029848f6",
  1025 => x"c087f8c0",
  1026 => x"c81ec0f4",
  1027 => x"87c70266",
  1028 => x"c048a6c4",
  1029 => x"c487c578",
  1030 => x"78c148a6",
  1031 => x"e74966c4",
  1032 => x"86c487d3",
  1033 => x"84c14d70",
  1034 => x"c14866c4",
  1035 => x"58a6c880",
  1036 => x"bfc0f0c2",
  1037 => x"c603ac49",
  1038 => x"059d7587",
  1039 => x"c087c8ff",
  1040 => x"029d754c",
  1041 => x"c087e0c3",
  1042 => x"c81ec0f4",
  1043 => x"87c70266",
  1044 => x"c048a6cc",
  1045 => x"cc87c578",
  1046 => x"78c148a6",
  1047 => x"e64966cc",
  1048 => x"86c487d3",
  1049 => x"98487e70",
  1050 => x"87e8c202",
  1051 => x"9781cb49",
  1052 => x"99d04969",
  1053 => x"87d6c102",
  1054 => x"4af6fec0",
  1055 => x"91cb4974",
  1056 => x"81dae0c1",
  1057 => x"81c87972",
  1058 => x"7451ffc3",
  1059 => x"c291de49",
  1060 => x"714dd4f0",
  1061 => x"97c1c285",
  1062 => x"49a5c17d",
  1063 => x"c251e0c0",
  1064 => x"bf97c6eb",
  1065 => x"c187d202",
  1066 => x"4ba5c284",
  1067 => x"4ac6ebc2",
  1068 => x"fffe49db",
  1069 => x"dbc187f1",
  1070 => x"49a5cd87",
  1071 => x"84c151c0",
  1072 => x"6e4ba5c2",
  1073 => x"fe49cb4a",
  1074 => x"c187dcff",
  1075 => x"fcc087c6",
  1076 => x"49744af2",
  1077 => x"e0c191cb",
  1078 => x"797281da",
  1079 => x"97c6ebc2",
  1080 => x"87d802bf",
  1081 => x"91de4974",
  1082 => x"f0c284c1",
  1083 => x"83714bd4",
  1084 => x"4ac6ebc2",
  1085 => x"fefe49dd",
  1086 => x"87d887ed",
  1087 => x"93de4b74",
  1088 => x"83d4f0c2",
  1089 => x"c049a3cb",
  1090 => x"7384c151",
  1091 => x"49cb4a6e",
  1092 => x"87d3fefe",
  1093 => x"c14866c4",
  1094 => x"58a6c880",
  1095 => x"c003acc7",
  1096 => x"056e87c5",
  1097 => x"7487e0fc",
  1098 => x"f68ef448",
  1099 => x"731e87ee",
  1100 => x"494b711e",
  1101 => x"e0c191cb",
  1102 => x"a1c881da",
  1103 => x"c6e0c14a",
  1104 => x"c9501248",
  1105 => x"f6c04aa1",
  1106 => x"501248ed",
  1107 => x"e0c181ca",
  1108 => x"501148c7",
  1109 => x"97c7e0c1",
  1110 => x"c01e49bf",
  1111 => x"87c3f749",
  1112 => x"48e8efc2",
  1113 => x"49c178de",
  1114 => x"2687e2d6",
  1115 => x"1e87f1f5",
  1116 => x"cb494a71",
  1117 => x"dae0c191",
  1118 => x"1181c881",
  1119 => x"ecefc248",
  1120 => x"c0f0c258",
  1121 => x"c178c048",
  1122 => x"87c1d649",
  1123 => x"c01e4f26",
  1124 => x"cbfbc049",
  1125 => x"1e4f2687",
  1126 => x"d2029971",
  1127 => x"efe1c187",
  1128 => x"f750c048",
  1129 => x"efc5c180",
  1130 => x"d3e0c140",
  1131 => x"c187ce78",
  1132 => x"c148ebe1",
  1133 => x"fc78cce0",
  1134 => x"cec6c180",
  1135 => x"0e4f2678",
  1136 => x"0e5c5b5e",
  1137 => x"cb4a4c71",
  1138 => x"dae0c192",
  1139 => x"49a2c882",
  1140 => x"974ba2c9",
  1141 => x"971e4b6b",
  1142 => x"ca1e4969",
  1143 => x"c0491282",
  1144 => x"c087c6e6",
  1145 => x"87e5d449",
  1146 => x"f8c04974",
  1147 => x"8ef887cd",
  1148 => x"1e87ebf3",
  1149 => x"4b711e73",
  1150 => x"87c3ff49",
  1151 => x"fefe4973",
  1152 => x"c049c087",
  1153 => x"f387d9f9",
  1154 => x"731e87d6",
  1155 => x"c64b711e",
  1156 => x"db024aa3",
  1157 => x"028ac187",
  1158 => x"028a87d6",
  1159 => x"8a87dac1",
  1160 => x"87fcc002",
  1161 => x"e1c0028a",
  1162 => x"cb028a87",
  1163 => x"87dbc187",
  1164 => x"fafc49c7",
  1165 => x"87dec187",
  1166 => x"bfc0f0c2",
  1167 => x"87cbc102",
  1168 => x"c288c148",
  1169 => x"c158c4f0",
  1170 => x"f0c287c1",
  1171 => x"c002bfc4",
  1172 => x"f0c287f9",
  1173 => x"c148bfc0",
  1174 => x"c4f0c280",
  1175 => x"87ebc058",
  1176 => x"bfc0f0c2",
  1177 => x"c289c649",
  1178 => x"c059c4f0",
  1179 => x"da03a9b7",
  1180 => x"c0f0c287",
  1181 => x"d278c048",
  1182 => x"c4f0c287",
  1183 => x"87cb02bf",
  1184 => x"bfc0f0c2",
  1185 => x"c280c648",
  1186 => x"c058c4f0",
  1187 => x"87fdd149",
  1188 => x"f5c04973",
  1189 => x"c7f187e5",
  1190 => x"5b5e0e87",
  1191 => x"ff0e5d5c",
  1192 => x"a6dc86d0",
  1193 => x"48a6c859",
  1194 => x"80c478c0",
  1195 => x"7866c4c1",
  1196 => x"78c180c4",
  1197 => x"78c180c4",
  1198 => x"48c4f0c2",
  1199 => x"efc278c1",
  1200 => x"de48bfe8",
  1201 => x"87cb05a8",
  1202 => x"7087d5f4",
  1203 => x"59a6cc49",
  1204 => x"e487f9cf",
  1205 => x"c5e587e3",
  1206 => x"87d2e487",
  1207 => x"fbc04c70",
  1208 => x"fbc102ac",
  1209 => x"0566d887",
  1210 => x"c187edc1",
  1211 => x"c44a66c0",
  1212 => x"727e6a82",
  1213 => x"c1dcc11e",
  1214 => x"4966c448",
  1215 => x"204aa1c8",
  1216 => x"05aa7141",
  1217 => x"511087f9",
  1218 => x"c0c14a26",
  1219 => x"c4c14866",
  1220 => x"496a78ee",
  1221 => x"517481c7",
  1222 => x"4966c0c1",
  1223 => x"51c181c8",
  1224 => x"4966c0c1",
  1225 => x"51c081c9",
  1226 => x"4966c0c1",
  1227 => x"51c081ca",
  1228 => x"1ed81ec1",
  1229 => x"81c8496a",
  1230 => x"c887f7e3",
  1231 => x"66c4c186",
  1232 => x"01a8c048",
  1233 => x"a6c887c7",
  1234 => x"ce78c148",
  1235 => x"66c4c187",
  1236 => x"d088c148",
  1237 => x"87c358a6",
  1238 => x"d087c3e3",
  1239 => x"78c248a6",
  1240 => x"cd029c74",
  1241 => x"66c887e2",
  1242 => x"66c8c148",
  1243 => x"d7cd03a8",
  1244 => x"48a6dc87",
  1245 => x"80e878c0",
  1246 => x"f1e178c0",
  1247 => x"c14c7087",
  1248 => x"c205acd0",
  1249 => x"66c487d7",
  1250 => x"87d5e47e",
  1251 => x"a6c84970",
  1252 => x"87dae159",
  1253 => x"ecc04c70",
  1254 => x"ebc105ac",
  1255 => x"4966c887",
  1256 => x"c0c191cb",
  1257 => x"a1c48166",
  1258 => x"c84d6a4a",
  1259 => x"66c44aa1",
  1260 => x"efc5c152",
  1261 => x"87f6e079",
  1262 => x"029c4c70",
  1263 => x"fbc087d8",
  1264 => x"87d202ac",
  1265 => x"e5e05574",
  1266 => x"9c4c7087",
  1267 => x"c087c702",
  1268 => x"ff05acfb",
  1269 => x"e0c087ee",
  1270 => x"55c1c255",
  1271 => x"d87d97c0",
  1272 => x"a96e4966",
  1273 => x"c887db05",
  1274 => x"66cc4866",
  1275 => x"87ca04a8",
  1276 => x"c14866c8",
  1277 => x"58a6cc80",
  1278 => x"66cc87c8",
  1279 => x"d088c148",
  1280 => x"dfff58a6",
  1281 => x"4c7087e8",
  1282 => x"05acd0c1",
  1283 => x"66d487c8",
  1284 => x"d880c148",
  1285 => x"d0c158a6",
  1286 => x"e9fd02ac",
  1287 => x"a6e0c087",
  1288 => x"7866d848",
  1289 => x"c04866c4",
  1290 => x"05a866e0",
  1291 => x"c087ebc9",
  1292 => x"c048a6e4",
  1293 => x"c0487478",
  1294 => x"7e7088fb",
  1295 => x"c9029848",
  1296 => x"cb4887ed",
  1297 => x"487e7088",
  1298 => x"cdc10298",
  1299 => x"88c94887",
  1300 => x"98487e70",
  1301 => x"87c1c402",
  1302 => x"7088c448",
  1303 => x"0298487e",
  1304 => x"c14887ce",
  1305 => x"487e7088",
  1306 => x"ecc30298",
  1307 => x"87e1c887",
  1308 => x"c048a6dc",
  1309 => x"ddff78f0",
  1310 => x"4c7087f4",
  1311 => x"02acecc0",
  1312 => x"c087c4c0",
  1313 => x"c05ca6e0",
  1314 => x"cd02acec",
  1315 => x"ddddff87",
  1316 => x"c04c7087",
  1317 => x"ff05acec",
  1318 => x"ecc087f3",
  1319 => x"c4c002ac",
  1320 => x"c9ddff87",
  1321 => x"ca1ec087",
  1322 => x"4966d01e",
  1323 => x"c8c191cb",
  1324 => x"80714866",
  1325 => x"c858a6cc",
  1326 => x"80c44866",
  1327 => x"cc58a6d0",
  1328 => x"ff49bf66",
  1329 => x"c187ebdd",
  1330 => x"d41ede1e",
  1331 => x"ff49bf66",
  1332 => x"d087dfdd",
  1333 => x"c0497086",
  1334 => x"ecc08909",
  1335 => x"e8c059a6",
  1336 => x"a8c04866",
  1337 => x"87eec006",
  1338 => x"4866e8c0",
  1339 => x"c003a8dd",
  1340 => x"66c487e4",
  1341 => x"e8c049bf",
  1342 => x"e0c08166",
  1343 => x"66e8c051",
  1344 => x"c481c149",
  1345 => x"c281bf66",
  1346 => x"e8c051c1",
  1347 => x"81c24966",
  1348 => x"81bf66c4",
  1349 => x"486e51c0",
  1350 => x"78eec4c1",
  1351 => x"81c8496e",
  1352 => x"6e5166d0",
  1353 => x"d481c949",
  1354 => x"496e5166",
  1355 => x"66dc81ca",
  1356 => x"4866d051",
  1357 => x"a6d480c1",
  1358 => x"4866c858",
  1359 => x"04a866cc",
  1360 => x"c887cbc0",
  1361 => x"80c14866",
  1362 => x"c558a6cc",
  1363 => x"66cc87e1",
  1364 => x"d088c148",
  1365 => x"d6c558a6",
  1366 => x"c4ddff87",
  1367 => x"c0497087",
  1368 => x"ff59a6ec",
  1369 => x"7087fadc",
  1370 => x"a6e0c049",
  1371 => x"4866dc59",
  1372 => x"05a8ecc0",
  1373 => x"dc87cac0",
  1374 => x"e8c048a6",
  1375 => x"c4c07866",
  1376 => x"e9d9ff87",
  1377 => x"4966c887",
  1378 => x"c0c191cb",
  1379 => x"80714866",
  1380 => x"c84a7e70",
  1381 => x"ca496e82",
  1382 => x"66e8c081",
  1383 => x"4966dc51",
  1384 => x"e8c081c1",
  1385 => x"48c18966",
  1386 => x"49703071",
  1387 => x"977189c1",
  1388 => x"f0f3c27a",
  1389 => x"e8c049bf",
  1390 => x"6a972966",
  1391 => x"9871484a",
  1392 => x"58a6f0c0",
  1393 => x"81c4496e",
  1394 => x"e0c04d69",
  1395 => x"66c44866",
  1396 => x"c8c002a8",
  1397 => x"48a6c487",
  1398 => x"c5c078c0",
  1399 => x"48a6c487",
  1400 => x"66c478c1",
  1401 => x"1ee0c01e",
  1402 => x"d9ff4975",
  1403 => x"86c887c4",
  1404 => x"b7c04c70",
  1405 => x"d4c106ac",
  1406 => x"c0857487",
  1407 => x"897449e0",
  1408 => x"dcc14b75",
  1409 => x"fe714aca",
  1410 => x"c287dcea",
  1411 => x"66e4c085",
  1412 => x"c080c148",
  1413 => x"c058a6e8",
  1414 => x"c14966ec",
  1415 => x"02a97081",
  1416 => x"c487c8c0",
  1417 => x"78c048a6",
  1418 => x"c487c5c0",
  1419 => x"78c148a6",
  1420 => x"c21e66c4",
  1421 => x"e0c049a4",
  1422 => x"70887148",
  1423 => x"49751e49",
  1424 => x"87eed7ff",
  1425 => x"b7c086c8",
  1426 => x"c0ff01a8",
  1427 => x"66e4c087",
  1428 => x"87d1c002",
  1429 => x"81c9496e",
  1430 => x"5166e4c0",
  1431 => x"c6c1486e",
  1432 => x"ccc078ff",
  1433 => x"c9496e87",
  1434 => x"6e51c281",
  1435 => x"f3c7c148",
  1436 => x"4866c878",
  1437 => x"04a866cc",
  1438 => x"c887cbc0",
  1439 => x"80c14866",
  1440 => x"c058a6cc",
  1441 => x"66cc87e9",
  1442 => x"d088c148",
  1443 => x"dec058a6",
  1444 => x"c9d6ff87",
  1445 => x"c04c7087",
  1446 => x"c6c187d5",
  1447 => x"c8c005ac",
  1448 => x"4866d087",
  1449 => x"a6d480c1",
  1450 => x"f1d5ff58",
  1451 => x"d44c7087",
  1452 => x"80c14866",
  1453 => x"7458a6d8",
  1454 => x"cbc0029c",
  1455 => x"4866c887",
  1456 => x"a866c8c1",
  1457 => x"87e9f204",
  1458 => x"87c9d5ff",
  1459 => x"c74866c8",
  1460 => x"e5c003a8",
  1461 => x"c4f0c287",
  1462 => x"c878c048",
  1463 => x"91cb4966",
  1464 => x"8166c0c1",
  1465 => x"6a4aa1c4",
  1466 => x"7952c04a",
  1467 => x"c14866c8",
  1468 => x"58a6cc80",
  1469 => x"ff04a8c7",
  1470 => x"d0ff87db",
  1471 => x"dbdfff8e",
  1472 => x"616f4c87",
  1473 => x"2e2a2064",
  1474 => x"203a0020",
  1475 => x"1e731e00",
  1476 => x"029b4b71",
  1477 => x"f0c287c6",
  1478 => x"78c048c0",
  1479 => x"f0c21ec7",
  1480 => x"1e49bfc0",
  1481 => x"1edae0c1",
  1482 => x"bfe8efc2",
  1483 => x"87e9ed49",
  1484 => x"efc286cc",
  1485 => x"e949bfe8",
  1486 => x"9b7387dd",
  1487 => x"c187c802",
  1488 => x"c049dae0",
  1489 => x"ff87c6e4",
  1490 => x"1e87d5de",
  1491 => x"4bc01e73",
  1492 => x"48c6e0c1",
  1493 => x"e1c150c0",
  1494 => x"ff49bffd",
  1495 => x"7087cfd9",
  1496 => x"87c40598",
  1497 => x"4beeddc1",
  1498 => x"ddff4873",
  1499 => x"4f5287f2",
  1500 => x"6f6c204d",
  1501 => x"6e696461",
  1502 => x"61662067",
  1503 => x"64656c69",
  1504 => x"dfc71e00",
  1505 => x"fe49c187",
  1506 => x"edfe87c3",
  1507 => x"987087ff",
  1508 => x"fe87cd02",
  1509 => x"7087d8f5",
  1510 => x"87c40298",
  1511 => x"87c24ac1",
  1512 => x"9a724ac0",
  1513 => x"c087ce05",
  1514 => x"d1dfc11e",
  1515 => x"d4efc049",
  1516 => x"fe86c487",
  1517 => x"c11ec087",
  1518 => x"c049dcdf",
  1519 => x"c087c6ef",
  1520 => x"87c7fe1e",
  1521 => x"eec04970",
  1522 => x"d6c387fb",
  1523 => x"268ef887",
  1524 => x"2044534f",
  1525 => x"6c696166",
  1526 => x"002e6465",
  1527 => x"746f6f42",
  1528 => x"2e676e69",
  1529 => x"1e002e2e",
  1530 => x"87dfe6c0",
  1531 => x"4f2687fa",
  1532 => x"c0f0c21e",
  1533 => x"c278c048",
  1534 => x"c048e8ef",
  1535 => x"87c1fe78",
  1536 => x"48c087e5",
  1537 => x"00004f26",
  1538 => x"00000001",
  1539 => x"78452080",
  1540 => x"80007469",
  1541 => x"63614220",
  1542 => x"0f32006b",
  1543 => x"2c140000",
  1544 => x"00000000",
  1545 => x"000f3200",
  1546 => x"002c3200",
  1547 => x"00000000",
  1548 => x"00000f32",
  1549 => x"00002c50",
  1550 => x"32000000",
  1551 => x"6e00000f",
  1552 => x"0000002c",
  1553 => x"0f320000",
  1554 => x"2c8c0000",
  1555 => x"00000000",
  1556 => x"000f3200",
  1557 => x"002caa00",
  1558 => x"00000000",
  1559 => x"00000f32",
  1560 => x"00002cc8",
  1561 => x"6f000000",
  1562 => x"00000011",
  1563 => x"00000000",
  1564 => x"120a0000",
  1565 => x"00000000",
  1566 => x"00000000",
  1567 => x"00188100",
  1568 => x"54455000",
  1569 => x"31303032",
  1570 => x"4d4f5220",
  1571 => x"f0fe1e00",
  1572 => x"cd78c048",
  1573 => x"26097909",
  1574 => x"fe1e1e4f",
  1575 => x"487ebff0",
  1576 => x"1e4f2626",
  1577 => x"c148f0fe",
  1578 => x"1e4f2678",
  1579 => x"c048f0fe",
  1580 => x"1e4f2678",
  1581 => x"52c04a71",
  1582 => x"0e4f2652",
  1583 => x"5d5c5b5e",
  1584 => x"7186f40e",
  1585 => x"7e6d974d",
  1586 => x"974ca5c1",
  1587 => x"a6c8486c",
  1588 => x"c4486e58",
  1589 => x"c505a866",
  1590 => x"c048ff87",
  1591 => x"caff87e6",
  1592 => x"49a5c287",
  1593 => x"714b6c97",
  1594 => x"6b974ba3",
  1595 => x"7e6c974b",
  1596 => x"80c1486e",
  1597 => x"c758a6c8",
  1598 => x"58a6cc98",
  1599 => x"fe7c9770",
  1600 => x"487387e1",
  1601 => x"4d268ef4",
  1602 => x"4b264c26",
  1603 => x"5e0e4f26",
  1604 => x"f40e5c5b",
  1605 => x"d84c7186",
  1606 => x"ffc34a66",
  1607 => x"4ba4c29a",
  1608 => x"73496c97",
  1609 => x"517249a1",
  1610 => x"6e7e6c97",
  1611 => x"c880c148",
  1612 => x"98c758a6",
  1613 => x"7058a6cc",
  1614 => x"ff8ef454",
  1615 => x"1e1e87ca",
  1616 => x"e087e8fd",
  1617 => x"c0494abf",
  1618 => x"0299c0e0",
  1619 => x"1e7287cb",
  1620 => x"49e6f3c2",
  1621 => x"c487f7fe",
  1622 => x"87fdfc86",
  1623 => x"c2fd7e70",
  1624 => x"4f262687",
  1625 => x"e6f3c21e",
  1626 => x"87c7fd49",
  1627 => x"49fee4c1",
  1628 => x"c387dafc",
  1629 => x"4f2687ee",
  1630 => x"5c5b5e0e",
  1631 => x"4d710e5d",
  1632 => x"49e6f3c2",
  1633 => x"7087f4fc",
  1634 => x"abb7c04b",
  1635 => x"87c2c304",
  1636 => x"05abf0c3",
  1637 => x"e9c187c9",
  1638 => x"78c148dc",
  1639 => x"c387e3c2",
  1640 => x"c905abe0",
  1641 => x"e0e9c187",
  1642 => x"c278c148",
  1643 => x"e9c187d4",
  1644 => x"c602bfe0",
  1645 => x"a3c0c287",
  1646 => x"7387c24c",
  1647 => x"dce9c14c",
  1648 => x"e0c002bf",
  1649 => x"c4497487",
  1650 => x"c19129b7",
  1651 => x"7481f3ea",
  1652 => x"c29acf4a",
  1653 => x"7248c192",
  1654 => x"ff4a7030",
  1655 => x"694872ba",
  1656 => x"db797098",
  1657 => x"c4497487",
  1658 => x"c19129b7",
  1659 => x"7481f3ea",
  1660 => x"c29acf4a",
  1661 => x"7248c392",
  1662 => x"484a7030",
  1663 => x"7970b069",
  1664 => x"c0059d75",
  1665 => x"d0ff87f0",
  1666 => x"78e1c848",
  1667 => x"c548d4ff",
  1668 => x"e0e9c178",
  1669 => x"87c302bf",
  1670 => x"c178e0c3",
  1671 => x"02bfdce9",
  1672 => x"d4ff87c6",
  1673 => x"78f0c348",
  1674 => x"7348d4ff",
  1675 => x"48d0ff78",
  1676 => x"c078e1c8",
  1677 => x"e9c178e0",
  1678 => x"78c048e0",
  1679 => x"48dce9c1",
  1680 => x"f3c278c0",
  1681 => x"f2f949e6",
  1682 => x"c04b7087",
  1683 => x"fc03abb7",
  1684 => x"48c087fe",
  1685 => x"4c264d26",
  1686 => x"4f264b26",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"724ac01e",
  1690 => x"c191c449",
  1691 => x"c081f3ea",
  1692 => x"d082c179",
  1693 => x"ee04aab7",
  1694 => x"0e4f2687",
  1695 => x"5d5c5b5e",
  1696 => x"f84d710e",
  1697 => x"4a7587e5",
  1698 => x"922ab7c4",
  1699 => x"82f3eac1",
  1700 => x"9ccf4c75",
  1701 => x"496a94c2",
  1702 => x"c32b744b",
  1703 => x"7448c29b",
  1704 => x"ff4c7030",
  1705 => x"714874bc",
  1706 => x"f77a7098",
  1707 => x"487387f5",
  1708 => x"0087e1fe",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000000",
  1717 => x"00000000",
  1718 => x"00000000",
  1719 => x"00000000",
  1720 => x"00000000",
  1721 => x"00000000",
  1722 => x"00000000",
  1723 => x"00000000",
  1724 => x"1e000000",
  1725 => x"c848d0ff",
  1726 => x"487178e1",
  1727 => x"7808d4ff",
  1728 => x"ff4866c4",
  1729 => x"267808d4",
  1730 => x"4a711e4f",
  1731 => x"1e4966c4",
  1732 => x"deff4972",
  1733 => x"48d0ff87",
  1734 => x"2678e0c0",
  1735 => x"731e4f26",
  1736 => x"c84b711e",
  1737 => x"731e4966",
  1738 => x"a2e0c14a",
  1739 => x"87d9ff49",
  1740 => x"2687c426",
  1741 => x"264c264d",
  1742 => x"1e4f264b",
  1743 => x"c34ad4ff",
  1744 => x"d0ff7aff",
  1745 => x"78e1c048",
  1746 => x"f3c27ade",
  1747 => x"497abff0",
  1748 => x"7028c848",
  1749 => x"d048717a",
  1750 => x"717a7028",
  1751 => x"7028d848",
  1752 => x"48d0ff7a",
  1753 => x"2678e0c0",
  1754 => x"5b5e0e4f",
  1755 => x"710e5d5c",
  1756 => x"f0f3c24c",
  1757 => x"74494dbf",
  1758 => x"d04b7129",
  1759 => x"83c19b66",
  1760 => x"abb766d4",
  1761 => x"c087c204",
  1762 => x"4966d04b",
  1763 => x"b9ff3174",
  1764 => x"4a739975",
  1765 => x"48723274",
  1766 => x"f3c2b071",
  1767 => x"dafe58f4",
  1768 => x"264d2687",
  1769 => x"264b264c",
  1770 => x"d0ff1e4f",
  1771 => x"78c9c848",
  1772 => x"d4ff4871",
  1773 => x"4f267808",
  1774 => x"494a711e",
  1775 => x"d0ff87eb",
  1776 => x"2678c848",
  1777 => x"1e731e4f",
  1778 => x"f4c24b71",
  1779 => x"c302bfc0",
  1780 => x"87ebc287",
  1781 => x"c848d0ff",
  1782 => x"497378c9",
  1783 => x"ffb1e0c0",
  1784 => x"787148d4",
  1785 => x"48f4f3c2",
  1786 => x"66c878c0",
  1787 => x"c387c502",
  1788 => x"87c249ff",
  1789 => x"f3c249c0",
  1790 => x"66cc59fc",
  1791 => x"c587c602",
  1792 => x"c44ad5d5",
  1793 => x"ffffcf87",
  1794 => x"c0f4c24a",
  1795 => x"c0f4c25a",
  1796 => x"c478c148",
  1797 => x"264d2687",
  1798 => x"264b264c",
  1799 => x"5b5e0e4f",
  1800 => x"710e5d5c",
  1801 => x"fcf3c24a",
  1802 => x"9a724cbf",
  1803 => x"4987cb02",
  1804 => x"eec191c8",
  1805 => x"83714bfb",
  1806 => x"f2c187c4",
  1807 => x"4dc04bfb",
  1808 => x"99744913",
  1809 => x"bff8f3c2",
  1810 => x"48d4ffb9",
  1811 => x"b7c17871",
  1812 => x"b7c8852c",
  1813 => x"87e804ad",
  1814 => x"bff4f3c2",
  1815 => x"c280c848",
  1816 => x"fe58f8f3",
  1817 => x"731e87ef",
  1818 => x"134b711e",
  1819 => x"cb029a4a",
  1820 => x"fe497287",
  1821 => x"4a1387e7",
  1822 => x"87f5059a",
  1823 => x"1e87dafe",
  1824 => x"bff4f3c2",
  1825 => x"f4f3c249",
  1826 => x"78a1c148",
  1827 => x"a9b7c0c4",
  1828 => x"ff87db03",
  1829 => x"f3c248d4",
  1830 => x"c278bff8",
  1831 => x"49bff4f3",
  1832 => x"48f4f3c2",
  1833 => x"c478a1c1",
  1834 => x"04a9b7c0",
  1835 => x"d0ff87e5",
  1836 => x"c278c848",
  1837 => x"c048c0f4",
  1838 => x"004f2678",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"5f5f0000",
  1842 => x"00000000",
  1843 => x"03000303",
  1844 => x"14000003",
  1845 => x"7f147f7f",
  1846 => x"0000147f",
  1847 => x"6b6b2e24",
  1848 => x"4c00123a",
  1849 => x"6c18366a",
  1850 => x"30003256",
  1851 => x"77594f7e",
  1852 => x"0040683a",
  1853 => x"03070400",
  1854 => x"00000000",
  1855 => x"633e1c00",
  1856 => x"00000041",
  1857 => x"3e634100",
  1858 => x"0800001c",
  1859 => x"1c1c3e2a",
  1860 => x"00082a3e",
  1861 => x"3e3e0808",
  1862 => x"00000808",
  1863 => x"60e08000",
  1864 => x"00000000",
  1865 => x"08080808",
  1866 => x"00000808",
  1867 => x"60600000",
  1868 => x"40000000",
  1869 => x"0c183060",
  1870 => x"00010306",
  1871 => x"4d597f3e",
  1872 => x"00003e7f",
  1873 => x"7f7f0604",
  1874 => x"00000000",
  1875 => x"59716342",
  1876 => x"0000464f",
  1877 => x"49496322",
  1878 => x"1800367f",
  1879 => x"7f13161c",
  1880 => x"0000107f",
  1881 => x"45456727",
  1882 => x"0000397d",
  1883 => x"494b7e3c",
  1884 => x"00003079",
  1885 => x"79710101",
  1886 => x"0000070f",
  1887 => x"49497f36",
  1888 => x"0000367f",
  1889 => x"69494f06",
  1890 => x"00001e3f",
  1891 => x"66660000",
  1892 => x"00000000",
  1893 => x"66e68000",
  1894 => x"00000000",
  1895 => x"14140808",
  1896 => x"00002222",
  1897 => x"14141414",
  1898 => x"00001414",
  1899 => x"14142222",
  1900 => x"00000808",
  1901 => x"59510302",
  1902 => x"3e00060f",
  1903 => x"555d417f",
  1904 => x"00001e1f",
  1905 => x"09097f7e",
  1906 => x"00007e7f",
  1907 => x"49497f7f",
  1908 => x"0000367f",
  1909 => x"41633e1c",
  1910 => x"00004141",
  1911 => x"63417f7f",
  1912 => x"00001c3e",
  1913 => x"49497f7f",
  1914 => x"00004141",
  1915 => x"09097f7f",
  1916 => x"00000101",
  1917 => x"49417f3e",
  1918 => x"00007a7b",
  1919 => x"08087f7f",
  1920 => x"00007f7f",
  1921 => x"7f7f4100",
  1922 => x"00000041",
  1923 => x"40406020",
  1924 => x"7f003f7f",
  1925 => x"361c087f",
  1926 => x"00004163",
  1927 => x"40407f7f",
  1928 => x"7f004040",
  1929 => x"060c067f",
  1930 => x"7f007f7f",
  1931 => x"180c067f",
  1932 => x"00007f7f",
  1933 => x"41417f3e",
  1934 => x"00003e7f",
  1935 => x"09097f7f",
  1936 => x"3e00060f",
  1937 => x"7f61417f",
  1938 => x"0000407e",
  1939 => x"19097f7f",
  1940 => x"0000667f",
  1941 => x"594d6f26",
  1942 => x"0000327b",
  1943 => x"7f7f0101",
  1944 => x"00000101",
  1945 => x"40407f3f",
  1946 => x"00003f7f",
  1947 => x"70703f0f",
  1948 => x"7f000f3f",
  1949 => x"3018307f",
  1950 => x"41007f7f",
  1951 => x"1c1c3663",
  1952 => x"01416336",
  1953 => x"7c7c0603",
  1954 => x"61010306",
  1955 => x"474d5971",
  1956 => x"00004143",
  1957 => x"417f7f00",
  1958 => x"01000041",
  1959 => x"180c0603",
  1960 => x"00406030",
  1961 => x"7f414100",
  1962 => x"0800007f",
  1963 => x"0603060c",
  1964 => x"8000080c",
  1965 => x"80808080",
  1966 => x"00008080",
  1967 => x"07030000",
  1968 => x"00000004",
  1969 => x"54547420",
  1970 => x"0000787c",
  1971 => x"44447f7f",
  1972 => x"0000387c",
  1973 => x"44447c38",
  1974 => x"00000044",
  1975 => x"44447c38",
  1976 => x"00007f7f",
  1977 => x"54547c38",
  1978 => x"0000185c",
  1979 => x"057f7e04",
  1980 => x"00000005",
  1981 => x"a4a4bc18",
  1982 => x"00007cfc",
  1983 => x"04047f7f",
  1984 => x"0000787c",
  1985 => x"7d3d0000",
  1986 => x"00000040",
  1987 => x"fd808080",
  1988 => x"0000007d",
  1989 => x"38107f7f",
  1990 => x"0000446c",
  1991 => x"7f3f0000",
  1992 => x"7c000040",
  1993 => x"0c180c7c",
  1994 => x"0000787c",
  1995 => x"04047c7c",
  1996 => x"0000787c",
  1997 => x"44447c38",
  1998 => x"0000387c",
  1999 => x"2424fcfc",
  2000 => x"0000183c",
  2001 => x"24243c18",
  2002 => x"0000fcfc",
  2003 => x"04047c7c",
  2004 => x"0000080c",
  2005 => x"54545c48",
  2006 => x"00002074",
  2007 => x"447f3f04",
  2008 => x"00000044",
  2009 => x"40407c3c",
  2010 => x"00007c7c",
  2011 => x"60603c1c",
  2012 => x"3c001c3c",
  2013 => x"6030607c",
  2014 => x"44003c7c",
  2015 => x"3810386c",
  2016 => x"0000446c",
  2017 => x"60e0bc1c",
  2018 => x"00001c3c",
  2019 => x"5c746444",
  2020 => x"0000444c",
  2021 => x"773e0808",
  2022 => x"00004141",
  2023 => x"7f7f0000",
  2024 => x"00000000",
  2025 => x"3e774141",
  2026 => x"02000808",
  2027 => x"02030101",
  2028 => x"7f000102",
  2029 => x"7f7f7f7f",
  2030 => x"08007f7f",
  2031 => x"3e1c1c08",
  2032 => x"7f7f7f3e",
  2033 => x"1c3e3e7f",
  2034 => x"0008081c",
  2035 => x"7c7c1810",
  2036 => x"00001018",
  2037 => x"7c7c3010",
  2038 => x"10001030",
  2039 => x"78606030",
  2040 => x"4200061e",
  2041 => x"3c183c66",
  2042 => x"78004266",
  2043 => x"c6c26a38",
  2044 => x"6000386c",
  2045 => x"00600000",
  2046 => x"0e006000",
  2047 => x"5d5c5b5e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
