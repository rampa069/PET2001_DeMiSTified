
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e0",x"f5",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e0",x"f5",x"c2"),
    14 => (x"48",x"d0",x"e2",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e5",x"de"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"9a",x"72",x"1e",x"73"),
    47 => (x"87",x"e7",x"c0",x"02"),
    48 => (x"4b",x"c1",x"48",x"c0"),
    49 => (x"d1",x"06",x"a9",x"72"),
    50 => (x"06",x"82",x"72",x"87"),
    51 => (x"83",x"73",x"87",x"c9"),
    52 => (x"f4",x"01",x"a9",x"72"),
    53 => (x"c1",x"87",x"c3",x"87"),
    54 => (x"a9",x"72",x"3a",x"b2"),
    55 => (x"80",x"73",x"89",x"03"),
    56 => (x"2b",x"2a",x"c1",x"07"),
    57 => (x"26",x"87",x"f3",x"05"),
    58 => (x"1e",x"4f",x"26",x"4b"),
    59 => (x"4d",x"c4",x"1e",x"75"),
    60 => (x"04",x"a1",x"b7",x"71"),
    61 => (x"81",x"c1",x"b9",x"ff"),
    62 => (x"72",x"07",x"bd",x"c3"),
    63 => (x"ff",x"04",x"a2",x"b7"),
    64 => (x"c1",x"82",x"c1",x"ba"),
    65 => (x"ee",x"fe",x"07",x"bd"),
    66 => (x"04",x"2d",x"c1",x"87"),
    67 => (x"80",x"c1",x"b8",x"ff"),
    68 => (x"ff",x"04",x"2d",x"07"),
    69 => (x"07",x"81",x"c1",x"b9"),
    70 => (x"4f",x"26",x"4d",x"26"),
    71 => (x"c4",x"4a",x"71",x"1e"),
    72 => (x"c1",x"48",x"49",x"66"),
    73 => (x"58",x"a6",x"c8",x"88"),
    74 => (x"d6",x"02",x"99",x"71"),
    75 => (x"48",x"d4",x"ff",x"87"),
    76 => (x"68",x"78",x"ff",x"c3"),
    77 => (x"49",x"66",x"c4",x"52"),
    78 => (x"c8",x"88",x"c1",x"48"),
    79 => (x"99",x"71",x"58",x"a6"),
    80 => (x"26",x"87",x"ea",x"05"),
    81 => (x"1e",x"73",x"1e",x"4f"),
    82 => (x"c3",x"4b",x"d4",x"ff"),
    83 => (x"4a",x"6b",x"7b",x"ff"),
    84 => (x"6b",x"7b",x"ff",x"c3"),
    85 => (x"72",x"32",x"c8",x"49"),
    86 => (x"7b",x"ff",x"c3",x"b1"),
    87 => (x"31",x"c8",x"4a",x"6b"),
    88 => (x"ff",x"c3",x"b2",x"71"),
    89 => (x"c8",x"49",x"6b",x"7b"),
    90 => (x"71",x"b1",x"72",x"32"),
    91 => (x"26",x"87",x"c4",x"48"),
    92 => (x"26",x"4c",x"26",x"4d"),
    93 => (x"0e",x"4f",x"26",x"4b"),
    94 => (x"5d",x"5c",x"5b",x"5e"),
    95 => (x"ff",x"4a",x"71",x"0e"),
    96 => (x"49",x"72",x"4c",x"d4"),
    97 => (x"71",x"99",x"ff",x"c3"),
    98 => (x"d0",x"e2",x"c2",x"7c"),
    99 => (x"87",x"c8",x"05",x"bf"),
   100 => (x"c9",x"48",x"66",x"d0"),
   101 => (x"58",x"a6",x"d4",x"30"),
   102 => (x"d8",x"49",x"66",x"d0"),
   103 => (x"99",x"ff",x"c3",x"29"),
   104 => (x"66",x"d0",x"7c",x"71"),
   105 => (x"c3",x"29",x"d0",x"49"),
   106 => (x"7c",x"71",x"99",x"ff"),
   107 => (x"c8",x"49",x"66",x"d0"),
   108 => (x"99",x"ff",x"c3",x"29"),
   109 => (x"66",x"d0",x"7c",x"71"),
   110 => (x"99",x"ff",x"c3",x"49"),
   111 => (x"49",x"72",x"7c",x"71"),
   112 => (x"ff",x"c3",x"29",x"d0"),
   113 => (x"6c",x"7c",x"71",x"99"),
   114 => (x"ff",x"f0",x"c9",x"4b"),
   115 => (x"ab",x"ff",x"c3",x"4d"),
   116 => (x"c3",x"87",x"d0",x"05"),
   117 => (x"4b",x"6c",x"7c",x"ff"),
   118 => (x"c6",x"02",x"8d",x"c1"),
   119 => (x"ab",x"ff",x"c3",x"87"),
   120 => (x"73",x"87",x"f0",x"02"),
   121 => (x"87",x"c7",x"fe",x"48"),
   122 => (x"ff",x"49",x"c0",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"c3",x"81",x"c1",x"78"),
   125 => (x"04",x"a9",x"b7",x"c8"),
   126 => (x"4f",x"26",x"87",x"f1"),
   127 => (x"e7",x"1e",x"73",x"1e"),
   128 => (x"df",x"f8",x"c4",x"87"),
   129 => (x"c0",x"1e",x"c0",x"4b"),
   130 => (x"f7",x"c1",x"f0",x"ff"),
   131 => (x"87",x"e7",x"fd",x"49"),
   132 => (x"a8",x"c1",x"86",x"c4"),
   133 => (x"87",x"ea",x"c0",x"05"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"c0",x"c1",x"78",x"ff"),
   136 => (x"c0",x"c0",x"c0",x"c0"),
   137 => (x"f0",x"e1",x"c0",x"1e"),
   138 => (x"fd",x"49",x"e9",x"c1"),
   139 => (x"86",x"c4",x"87",x"c9"),
   140 => (x"ca",x"05",x"98",x"70"),
   141 => (x"48",x"d4",x"ff",x"87"),
   142 => (x"c1",x"78",x"ff",x"c3"),
   143 => (x"fe",x"87",x"cb",x"48"),
   144 => (x"8b",x"c1",x"87",x"e6"),
   145 => (x"87",x"fd",x"fe",x"05"),
   146 => (x"e6",x"fc",x"48",x"c0"),
   147 => (x"1e",x"73",x"1e",x"87"),
   148 => (x"c3",x"48",x"d4",x"ff"),
   149 => (x"4b",x"d3",x"78",x"ff"),
   150 => (x"ff",x"c0",x"1e",x"c0"),
   151 => (x"49",x"c1",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d4",x"fc"),
   153 => (x"05",x"98",x"70",x"86"),
   154 => (x"d4",x"ff",x"87",x"ca"),
   155 => (x"78",x"ff",x"c3",x"48"),
   156 => (x"87",x"cb",x"48",x"c1"),
   157 => (x"c1",x"87",x"f1",x"fd"),
   158 => (x"db",x"ff",x"05",x"8b"),
   159 => (x"fb",x"48",x"c0",x"87"),
   160 => (x"5e",x"0e",x"87",x"f1"),
   161 => (x"ff",x"0e",x"5c",x"5b"),
   162 => (x"db",x"fd",x"4c",x"d4"),
   163 => (x"1e",x"ea",x"c6",x"87"),
   164 => (x"c1",x"f0",x"e1",x"c0"),
   165 => (x"de",x"fb",x"49",x"c8"),
   166 => (x"c1",x"86",x"c4",x"87"),
   167 => (x"87",x"c8",x"02",x"a8"),
   168 => (x"c0",x"87",x"ea",x"fe"),
   169 => (x"87",x"e2",x"c1",x"48"),
   170 => (x"70",x"87",x"da",x"fa"),
   171 => (x"ff",x"ff",x"cf",x"49"),
   172 => (x"a9",x"ea",x"c6",x"99"),
   173 => (x"fe",x"87",x"c8",x"02"),
   174 => (x"48",x"c0",x"87",x"d3"),
   175 => (x"c3",x"87",x"cb",x"c1"),
   176 => (x"f1",x"c0",x"7c",x"ff"),
   177 => (x"87",x"f4",x"fc",x"4b"),
   178 => (x"c0",x"02",x"98",x"70"),
   179 => (x"1e",x"c0",x"87",x"eb"),
   180 => (x"c1",x"f0",x"ff",x"c0"),
   181 => (x"de",x"fa",x"49",x"fa"),
   182 => (x"70",x"86",x"c4",x"87"),
   183 => (x"87",x"d9",x"05",x"98"),
   184 => (x"6c",x"7c",x"ff",x"c3"),
   185 => (x"7c",x"ff",x"c3",x"49"),
   186 => (x"c1",x"7c",x"7c",x"7c"),
   187 => (x"c4",x"02",x"99",x"c0"),
   188 => (x"d5",x"48",x"c1",x"87"),
   189 => (x"d1",x"48",x"c0",x"87"),
   190 => (x"05",x"ab",x"c2",x"87"),
   191 => (x"48",x"c0",x"87",x"c4"),
   192 => (x"8b",x"c1",x"87",x"c8"),
   193 => (x"87",x"fd",x"fe",x"05"),
   194 => (x"e4",x"f9",x"48",x"c0"),
   195 => (x"1e",x"73",x"1e",x"87"),
   196 => (x"48",x"d0",x"e2",x"c2"),
   197 => (x"4b",x"c7",x"78",x"c1"),
   198 => (x"c2",x"48",x"d0",x"ff"),
   199 => (x"87",x"c8",x"fb",x"78"),
   200 => (x"c3",x"48",x"d0",x"ff"),
   201 => (x"c0",x"1e",x"c0",x"78"),
   202 => (x"c0",x"c1",x"d0",x"e5"),
   203 => (x"87",x"c7",x"f9",x"49"),
   204 => (x"a8",x"c1",x"86",x"c4"),
   205 => (x"4b",x"87",x"c1",x"05"),
   206 => (x"c5",x"05",x"ab",x"c2"),
   207 => (x"c0",x"48",x"c0",x"87"),
   208 => (x"8b",x"c1",x"87",x"f9"),
   209 => (x"87",x"d0",x"ff",x"05"),
   210 => (x"c2",x"87",x"f7",x"fc"),
   211 => (x"70",x"58",x"d4",x"e2"),
   212 => (x"87",x"cd",x"05",x"98"),
   213 => (x"ff",x"c0",x"1e",x"c1"),
   214 => (x"49",x"d0",x"c1",x"f0"),
   215 => (x"c4",x"87",x"d8",x"f8"),
   216 => (x"48",x"d4",x"ff",x"86"),
   217 => (x"c2",x"78",x"ff",x"c3"),
   218 => (x"e2",x"c2",x"87",x"fc"),
   219 => (x"d0",x"ff",x"58",x"d8"),
   220 => (x"ff",x"78",x"c2",x"48"),
   221 => (x"ff",x"c3",x"48",x"d4"),
   222 => (x"f7",x"48",x"c1",x"78"),
   223 => (x"5e",x"0e",x"87",x"f5"),
   224 => (x"0e",x"5d",x"5c",x"5b"),
   225 => (x"4c",x"c0",x"4b",x"71"),
   226 => (x"df",x"cd",x"ee",x"c5"),
   227 => (x"48",x"d4",x"ff",x"4a"),
   228 => (x"68",x"78",x"ff",x"c3"),
   229 => (x"a9",x"fe",x"c3",x"49"),
   230 => (x"87",x"fd",x"c0",x"05"),
   231 => (x"9b",x"73",x"4d",x"70"),
   232 => (x"d0",x"87",x"cc",x"02"),
   233 => (x"49",x"73",x"1e",x"66"),
   234 => (x"c4",x"87",x"f1",x"f5"),
   235 => (x"ff",x"87",x"d6",x"86"),
   236 => (x"d1",x"c4",x"48",x"d0"),
   237 => (x"7d",x"ff",x"c3",x"78"),
   238 => (x"c1",x"48",x"66",x"d0"),
   239 => (x"58",x"a6",x"d4",x"88"),
   240 => (x"f0",x"05",x"98",x"70"),
   241 => (x"48",x"d4",x"ff",x"87"),
   242 => (x"78",x"78",x"ff",x"c3"),
   243 => (x"c5",x"05",x"9b",x"73"),
   244 => (x"48",x"d0",x"ff",x"87"),
   245 => (x"4a",x"c1",x"78",x"d0"),
   246 => (x"05",x"8a",x"c1",x"4c"),
   247 => (x"74",x"87",x"ee",x"fe"),
   248 => (x"87",x"cb",x"f6",x"48"),
   249 => (x"71",x"1e",x"73",x"1e"),
   250 => (x"ff",x"4b",x"c0",x"4a"),
   251 => (x"ff",x"c3",x"48",x"d4"),
   252 => (x"48",x"d0",x"ff",x"78"),
   253 => (x"ff",x"78",x"c3",x"c4"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"c0",x"1e",x"72",x"78"),
   256 => (x"d1",x"c1",x"f0",x"ff"),
   257 => (x"87",x"ef",x"f5",x"49"),
   258 => (x"98",x"70",x"86",x"c4"),
   259 => (x"c8",x"87",x"d2",x"05"),
   260 => (x"66",x"cc",x"1e",x"c0"),
   261 => (x"87",x"e6",x"fd",x"49"),
   262 => (x"4b",x"70",x"86",x"c4"),
   263 => (x"c2",x"48",x"d0",x"ff"),
   264 => (x"f5",x"48",x"73",x"78"),
   265 => (x"5e",x"0e",x"87",x"cd"),
   266 => (x"0e",x"5d",x"5c",x"5b"),
   267 => (x"ff",x"c0",x"1e",x"c0"),
   268 => (x"49",x"c9",x"c1",x"f0"),
   269 => (x"d2",x"87",x"c0",x"f5"),
   270 => (x"d8",x"e2",x"c2",x"1e"),
   271 => (x"87",x"fe",x"fc",x"49"),
   272 => (x"4c",x"c0",x"86",x"c8"),
   273 => (x"b7",x"d2",x"84",x"c1"),
   274 => (x"87",x"f8",x"04",x"ac"),
   275 => (x"97",x"d8",x"e2",x"c2"),
   276 => (x"c0",x"c3",x"49",x"bf"),
   277 => (x"a9",x"c0",x"c1",x"99"),
   278 => (x"87",x"e7",x"c0",x"05"),
   279 => (x"97",x"df",x"e2",x"c2"),
   280 => (x"31",x"d0",x"49",x"bf"),
   281 => (x"97",x"e0",x"e2",x"c2"),
   282 => (x"32",x"c8",x"4a",x"bf"),
   283 => (x"e2",x"c2",x"b1",x"72"),
   284 => (x"4a",x"bf",x"97",x"e1"),
   285 => (x"cf",x"4c",x"71",x"b1"),
   286 => (x"9c",x"ff",x"ff",x"ff"),
   287 => (x"34",x"ca",x"84",x"c1"),
   288 => (x"c2",x"87",x"e7",x"c1"),
   289 => (x"bf",x"97",x"e1",x"e2"),
   290 => (x"c6",x"31",x"c1",x"49"),
   291 => (x"e2",x"e2",x"c2",x"99"),
   292 => (x"c7",x"4a",x"bf",x"97"),
   293 => (x"b1",x"72",x"2a",x"b7"),
   294 => (x"97",x"dd",x"e2",x"c2"),
   295 => (x"cf",x"4d",x"4a",x"bf"),
   296 => (x"de",x"e2",x"c2",x"9d"),
   297 => (x"c3",x"4a",x"bf",x"97"),
   298 => (x"c2",x"32",x"ca",x"9a"),
   299 => (x"bf",x"97",x"df",x"e2"),
   300 => (x"73",x"33",x"c2",x"4b"),
   301 => (x"e0",x"e2",x"c2",x"b2"),
   302 => (x"c3",x"4b",x"bf",x"97"),
   303 => (x"b7",x"c6",x"9b",x"c0"),
   304 => (x"c2",x"b2",x"73",x"2b"),
   305 => (x"71",x"48",x"c1",x"81"),
   306 => (x"c1",x"49",x"70",x"30"),
   307 => (x"70",x"30",x"75",x"48"),
   308 => (x"c1",x"4c",x"72",x"4d"),
   309 => (x"c8",x"94",x"71",x"84"),
   310 => (x"06",x"ad",x"b7",x"c0"),
   311 => (x"34",x"c1",x"87",x"cc"),
   312 => (x"c0",x"c8",x"2d",x"b7"),
   313 => (x"ff",x"01",x"ad",x"b7"),
   314 => (x"48",x"74",x"87",x"f4"),
   315 => (x"0e",x"87",x"c0",x"f2"),
   316 => (x"5d",x"5c",x"5b",x"5e"),
   317 => (x"c2",x"86",x"f8",x"0e"),
   318 => (x"c0",x"48",x"fe",x"ea"),
   319 => (x"f6",x"e2",x"c2",x"78"),
   320 => (x"fb",x"49",x"c0",x"1e"),
   321 => (x"86",x"c4",x"87",x"de"),
   322 => (x"c5",x"05",x"98",x"70"),
   323 => (x"c9",x"48",x"c0",x"87"),
   324 => (x"4d",x"c0",x"87",x"ce"),
   325 => (x"ef",x"c0",x"7e",x"c1"),
   326 => (x"c2",x"49",x"bf",x"d8"),
   327 => (x"71",x"4a",x"ec",x"e3"),
   328 => (x"c4",x"ed",x"4b",x"c8"),
   329 => (x"05",x"98",x"70",x"87"),
   330 => (x"7e",x"c0",x"87",x"c2"),
   331 => (x"bf",x"d4",x"ef",x"c0"),
   332 => (x"c8",x"e4",x"c2",x"49"),
   333 => (x"4b",x"c8",x"71",x"4a"),
   334 => (x"70",x"87",x"ee",x"ec"),
   335 => (x"87",x"c2",x"05",x"98"),
   336 => (x"02",x"6e",x"7e",x"c0"),
   337 => (x"c2",x"87",x"fd",x"c0"),
   338 => (x"4d",x"bf",x"fc",x"e9"),
   339 => (x"9f",x"f4",x"ea",x"c2"),
   340 => (x"c5",x"48",x"7e",x"bf"),
   341 => (x"05",x"a8",x"ea",x"d6"),
   342 => (x"e9",x"c2",x"87",x"c7"),
   343 => (x"ce",x"4d",x"bf",x"fc"),
   344 => (x"ca",x"48",x"6e",x"87"),
   345 => (x"02",x"a8",x"d5",x"e9"),
   346 => (x"48",x"c0",x"87",x"c5"),
   347 => (x"c2",x"87",x"f1",x"c7"),
   348 => (x"75",x"1e",x"f6",x"e2"),
   349 => (x"87",x"ec",x"f9",x"49"),
   350 => (x"98",x"70",x"86",x"c4"),
   351 => (x"c0",x"87",x"c5",x"05"),
   352 => (x"87",x"dc",x"c7",x"48"),
   353 => (x"bf",x"d4",x"ef",x"c0"),
   354 => (x"c8",x"e4",x"c2",x"49"),
   355 => (x"4b",x"c8",x"71",x"4a"),
   356 => (x"70",x"87",x"d6",x"eb"),
   357 => (x"87",x"c8",x"05",x"98"),
   358 => (x"48",x"fe",x"ea",x"c2"),
   359 => (x"87",x"da",x"78",x"c1"),
   360 => (x"bf",x"d8",x"ef",x"c0"),
   361 => (x"ec",x"e3",x"c2",x"49"),
   362 => (x"4b",x"c8",x"71",x"4a"),
   363 => (x"70",x"87",x"fa",x"ea"),
   364 => (x"c5",x"c0",x"02",x"98"),
   365 => (x"c6",x"48",x"c0",x"87"),
   366 => (x"ea",x"c2",x"87",x"e6"),
   367 => (x"49",x"bf",x"97",x"f4"),
   368 => (x"05",x"a9",x"d5",x"c1"),
   369 => (x"c2",x"87",x"cd",x"c0"),
   370 => (x"bf",x"97",x"f5",x"ea"),
   371 => (x"a9",x"ea",x"c2",x"49"),
   372 => (x"87",x"c5",x"c0",x"02"),
   373 => (x"c7",x"c6",x"48",x"c0"),
   374 => (x"f6",x"e2",x"c2",x"87"),
   375 => (x"48",x"7e",x"bf",x"97"),
   376 => (x"02",x"a8",x"e9",x"c3"),
   377 => (x"6e",x"87",x"ce",x"c0"),
   378 => (x"a8",x"eb",x"c3",x"48"),
   379 => (x"87",x"c5",x"c0",x"02"),
   380 => (x"eb",x"c5",x"48",x"c0"),
   381 => (x"c1",x"e3",x"c2",x"87"),
   382 => (x"99",x"49",x"bf",x"97"),
   383 => (x"87",x"cc",x"c0",x"05"),
   384 => (x"97",x"c2",x"e3",x"c2"),
   385 => (x"a9",x"c2",x"49",x"bf"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"cf",x"c5",x"48",x"c0"),
   388 => (x"c3",x"e3",x"c2",x"87"),
   389 => (x"c2",x"48",x"bf",x"97"),
   390 => (x"70",x"58",x"fa",x"ea"),
   391 => (x"88",x"c1",x"48",x"4c"),
   392 => (x"58",x"fe",x"ea",x"c2"),
   393 => (x"97",x"c4",x"e3",x"c2"),
   394 => (x"81",x"75",x"49",x"bf"),
   395 => (x"97",x"c5",x"e3",x"c2"),
   396 => (x"32",x"c8",x"4a",x"bf"),
   397 => (x"c2",x"7e",x"a1",x"72"),
   398 => (x"6e",x"48",x"cb",x"ef"),
   399 => (x"c6",x"e3",x"c2",x"78"),
   400 => (x"c8",x"48",x"bf",x"97"),
   401 => (x"ea",x"c2",x"58",x"a6"),
   402 => (x"c2",x"02",x"bf",x"fe"),
   403 => (x"ef",x"c0",x"87",x"d4"),
   404 => (x"c2",x"49",x"bf",x"d4"),
   405 => (x"71",x"4a",x"c8",x"e4"),
   406 => (x"cc",x"e8",x"4b",x"c8"),
   407 => (x"02",x"98",x"70",x"87"),
   408 => (x"c0",x"87",x"c5",x"c0"),
   409 => (x"87",x"f8",x"c3",x"48"),
   410 => (x"bf",x"f6",x"ea",x"c2"),
   411 => (x"df",x"ef",x"c2",x"4c"),
   412 => (x"db",x"e3",x"c2",x"5c"),
   413 => (x"c8",x"49",x"bf",x"97"),
   414 => (x"da",x"e3",x"c2",x"31"),
   415 => (x"a1",x"4a",x"bf",x"97"),
   416 => (x"dc",x"e3",x"c2",x"49"),
   417 => (x"d0",x"4a",x"bf",x"97"),
   418 => (x"49",x"a1",x"72",x"32"),
   419 => (x"97",x"dd",x"e3",x"c2"),
   420 => (x"32",x"d8",x"4a",x"bf"),
   421 => (x"c4",x"49",x"a1",x"72"),
   422 => (x"ef",x"c2",x"91",x"66"),
   423 => (x"c2",x"81",x"bf",x"cb"),
   424 => (x"c2",x"59",x"d3",x"ef"),
   425 => (x"bf",x"97",x"e3",x"e3"),
   426 => (x"c2",x"32",x"c8",x"4a"),
   427 => (x"bf",x"97",x"e2",x"e3"),
   428 => (x"c2",x"4a",x"a2",x"4b"),
   429 => (x"bf",x"97",x"e4",x"e3"),
   430 => (x"73",x"33",x"d0",x"4b"),
   431 => (x"e3",x"c2",x"4a",x"a2"),
   432 => (x"4b",x"bf",x"97",x"e5"),
   433 => (x"33",x"d8",x"9b",x"cf"),
   434 => (x"c2",x"4a",x"a2",x"73"),
   435 => (x"c2",x"5a",x"d7",x"ef"),
   436 => (x"4a",x"bf",x"d3",x"ef"),
   437 => (x"92",x"74",x"8a",x"c2"),
   438 => (x"48",x"d7",x"ef",x"c2"),
   439 => (x"c1",x"78",x"a1",x"72"),
   440 => (x"e3",x"c2",x"87",x"ca"),
   441 => (x"49",x"bf",x"97",x"c8"),
   442 => (x"e3",x"c2",x"31",x"c8"),
   443 => (x"4a",x"bf",x"97",x"c7"),
   444 => (x"eb",x"c2",x"49",x"a1"),
   445 => (x"eb",x"c2",x"59",x"c6"),
   446 => (x"c5",x"49",x"bf",x"c2"),
   447 => (x"81",x"ff",x"c7",x"31"),
   448 => (x"ef",x"c2",x"29",x"c9"),
   449 => (x"e3",x"c2",x"59",x"df"),
   450 => (x"4a",x"bf",x"97",x"cd"),
   451 => (x"e3",x"c2",x"32",x"c8"),
   452 => (x"4b",x"bf",x"97",x"cc"),
   453 => (x"66",x"c4",x"4a",x"a2"),
   454 => (x"c2",x"82",x"6e",x"92"),
   455 => (x"c2",x"5a",x"db",x"ef"),
   456 => (x"c0",x"48",x"d3",x"ef"),
   457 => (x"cf",x"ef",x"c2",x"78"),
   458 => (x"78",x"a1",x"72",x"48"),
   459 => (x"48",x"df",x"ef",x"c2"),
   460 => (x"bf",x"d3",x"ef",x"c2"),
   461 => (x"e3",x"ef",x"c2",x"78"),
   462 => (x"d7",x"ef",x"c2",x"48"),
   463 => (x"ea",x"c2",x"78",x"bf"),
   464 => (x"c0",x"02",x"bf",x"fe"),
   465 => (x"48",x"74",x"87",x"c9"),
   466 => (x"7e",x"70",x"30",x"c4"),
   467 => (x"c2",x"87",x"c9",x"c0"),
   468 => (x"48",x"bf",x"db",x"ef"),
   469 => (x"7e",x"70",x"30",x"c4"),
   470 => (x"48",x"c2",x"eb",x"c2"),
   471 => (x"48",x"c1",x"78",x"6e"),
   472 => (x"4d",x"26",x"8e",x"f8"),
   473 => (x"4b",x"26",x"4c",x"26"),
   474 => (x"5e",x"0e",x"4f",x"26"),
   475 => (x"0e",x"5d",x"5c",x"5b"),
   476 => (x"ea",x"c2",x"4a",x"71"),
   477 => (x"cb",x"02",x"bf",x"fe"),
   478 => (x"c7",x"4b",x"72",x"87"),
   479 => (x"c1",x"4c",x"72",x"2b"),
   480 => (x"87",x"c9",x"9c",x"ff"),
   481 => (x"2b",x"c8",x"4b",x"72"),
   482 => (x"ff",x"c3",x"4c",x"72"),
   483 => (x"cb",x"ef",x"c2",x"9c"),
   484 => (x"ef",x"c0",x"83",x"bf"),
   485 => (x"02",x"ab",x"bf",x"d0"),
   486 => (x"ef",x"c0",x"87",x"d9"),
   487 => (x"e2",x"c2",x"5b",x"d4"),
   488 => (x"49",x"73",x"1e",x"f6"),
   489 => (x"c4",x"87",x"fd",x"f0"),
   490 => (x"05",x"98",x"70",x"86"),
   491 => (x"48",x"c0",x"87",x"c5"),
   492 => (x"c2",x"87",x"e6",x"c0"),
   493 => (x"02",x"bf",x"fe",x"ea"),
   494 => (x"49",x"74",x"87",x"d2"),
   495 => (x"e2",x"c2",x"91",x"c4"),
   496 => (x"4d",x"69",x"81",x"f6"),
   497 => (x"ff",x"ff",x"ff",x"cf"),
   498 => (x"87",x"cb",x"9d",x"ff"),
   499 => (x"91",x"c2",x"49",x"74"),
   500 => (x"81",x"f6",x"e2",x"c2"),
   501 => (x"75",x"4d",x"69",x"9f"),
   502 => (x"87",x"c6",x"fe",x"48"),
   503 => (x"5c",x"5b",x"5e",x"0e"),
   504 => (x"86",x"f8",x"0e",x"5d"),
   505 => (x"05",x"9c",x"4c",x"71"),
   506 => (x"48",x"c0",x"87",x"c5"),
   507 => (x"c8",x"87",x"c2",x"c3"),
   508 => (x"48",x"6e",x"7e",x"a4"),
   509 => (x"66",x"d8",x"78",x"c0"),
   510 => (x"d8",x"87",x"c7",x"02"),
   511 => (x"05",x"bf",x"97",x"66"),
   512 => (x"48",x"c0",x"87",x"c5"),
   513 => (x"c0",x"87",x"ea",x"c2"),
   514 => (x"49",x"49",x"c1",x"1e"),
   515 => (x"c4",x"87",x"e6",x"c7"),
   516 => (x"9d",x"4d",x"70",x"86"),
   517 => (x"87",x"c2",x"c1",x"02"),
   518 => (x"4a",x"c6",x"eb",x"c2"),
   519 => (x"e0",x"49",x"66",x"d8"),
   520 => (x"98",x"70",x"87",x"ec"),
   521 => (x"87",x"f2",x"c0",x"02"),
   522 => (x"66",x"d8",x"4a",x"75"),
   523 => (x"e1",x"4b",x"cb",x"49"),
   524 => (x"98",x"70",x"87",x"d1"),
   525 => (x"87",x"e2",x"c0",x"02"),
   526 => (x"9d",x"75",x"1e",x"c0"),
   527 => (x"c8",x"87",x"c7",x"02"),
   528 => (x"78",x"c0",x"48",x"a6"),
   529 => (x"a6",x"c8",x"87",x"c5"),
   530 => (x"c8",x"78",x"c1",x"48"),
   531 => (x"e4",x"c6",x"49",x"66"),
   532 => (x"70",x"86",x"c4",x"87"),
   533 => (x"fe",x"05",x"9d",x"4d"),
   534 => (x"9d",x"75",x"87",x"fe"),
   535 => (x"87",x"cf",x"c1",x"02"),
   536 => (x"6e",x"49",x"a5",x"dc"),
   537 => (x"da",x"78",x"69",x"48"),
   538 => (x"a6",x"c4",x"49",x"a5"),
   539 => (x"78",x"a4",x"c4",x"48"),
   540 => (x"c4",x"48",x"69",x"9f"),
   541 => (x"c2",x"78",x"08",x"66"),
   542 => (x"02",x"bf",x"fe",x"ea"),
   543 => (x"a5",x"d4",x"87",x"d2"),
   544 => (x"49",x"69",x"9f",x"49"),
   545 => (x"99",x"ff",x"ff",x"c0"),
   546 => (x"30",x"d0",x"48",x"71"),
   547 => (x"87",x"c2",x"7e",x"70"),
   548 => (x"49",x"6e",x"7e",x"c0"),
   549 => (x"bf",x"66",x"c4",x"48"),
   550 => (x"08",x"66",x"c4",x"80"),
   551 => (x"cc",x"7c",x"c0",x"78"),
   552 => (x"66",x"c4",x"49",x"a4"),
   553 => (x"a4",x"d0",x"79",x"bf"),
   554 => (x"c1",x"79",x"c0",x"49"),
   555 => (x"c0",x"87",x"c2",x"48"),
   556 => (x"fa",x"8e",x"f8",x"48"),
   557 => (x"5e",x"0e",x"87",x"ec"),
   558 => (x"0e",x"5d",x"5c",x"5b"),
   559 => (x"02",x"9c",x"4c",x"71"),
   560 => (x"c8",x"87",x"ca",x"c1"),
   561 => (x"02",x"69",x"49",x"a4"),
   562 => (x"d0",x"87",x"c2",x"c1"),
   563 => (x"49",x"6c",x"4a",x"66"),
   564 => (x"5a",x"a6",x"d4",x"82"),
   565 => (x"b9",x"4d",x"66",x"d0"),
   566 => (x"bf",x"fa",x"ea",x"c2"),
   567 => (x"72",x"ba",x"ff",x"4a"),
   568 => (x"02",x"99",x"71",x"99"),
   569 => (x"c4",x"87",x"e4",x"c0"),
   570 => (x"49",x"6b",x"4b",x"a4"),
   571 => (x"70",x"87",x"fb",x"f9"),
   572 => (x"f6",x"ea",x"c2",x"7b"),
   573 => (x"81",x"6c",x"49",x"bf"),
   574 => (x"b9",x"75",x"7c",x"71"),
   575 => (x"bf",x"fa",x"ea",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"05",x"99",x"71",x"99"),
   578 => (x"75",x"87",x"dc",x"ff"),
   579 => (x"87",x"d2",x"f9",x"7c"),
   580 => (x"71",x"1e",x"73",x"1e"),
   581 => (x"c7",x"02",x"9b",x"4b"),
   582 => (x"49",x"a3",x"c8",x"87"),
   583 => (x"87",x"c5",x"05",x"69"),
   584 => (x"f7",x"c0",x"48",x"c0"),
   585 => (x"cf",x"ef",x"c2",x"87"),
   586 => (x"a3",x"c4",x"4a",x"bf"),
   587 => (x"c2",x"49",x"69",x"49"),
   588 => (x"f6",x"ea",x"c2",x"89"),
   589 => (x"a2",x"71",x"91",x"bf"),
   590 => (x"fa",x"ea",x"c2",x"4a"),
   591 => (x"99",x"6b",x"49",x"bf"),
   592 => (x"c0",x"4a",x"a2",x"71"),
   593 => (x"c8",x"5a",x"d4",x"ef"),
   594 => (x"49",x"72",x"1e",x"66"),
   595 => (x"c4",x"87",x"d5",x"ea"),
   596 => (x"05",x"98",x"70",x"86"),
   597 => (x"48",x"c0",x"87",x"c4"),
   598 => (x"48",x"c1",x"87",x"c2"),
   599 => (x"1e",x"87",x"c7",x"f8"),
   600 => (x"4b",x"71",x"1e",x"73"),
   601 => (x"e4",x"c0",x"02",x"9b"),
   602 => (x"e3",x"ef",x"c2",x"87"),
   603 => (x"c2",x"4a",x"73",x"5b"),
   604 => (x"f6",x"ea",x"c2",x"8a"),
   605 => (x"c2",x"92",x"49",x"bf"),
   606 => (x"48",x"bf",x"cf",x"ef"),
   607 => (x"ef",x"c2",x"80",x"72"),
   608 => (x"48",x"71",x"58",x"e7"),
   609 => (x"eb",x"c2",x"30",x"c4"),
   610 => (x"ed",x"c0",x"58",x"c6"),
   611 => (x"df",x"ef",x"c2",x"87"),
   612 => (x"d3",x"ef",x"c2",x"48"),
   613 => (x"ef",x"c2",x"78",x"bf"),
   614 => (x"ef",x"c2",x"48",x"e3"),
   615 => (x"c2",x"78",x"bf",x"d7"),
   616 => (x"02",x"bf",x"fe",x"ea"),
   617 => (x"ea",x"c2",x"87",x"c9"),
   618 => (x"c4",x"49",x"bf",x"f6"),
   619 => (x"c2",x"87",x"c7",x"31"),
   620 => (x"49",x"bf",x"db",x"ef"),
   621 => (x"eb",x"c2",x"31",x"c4"),
   622 => (x"e9",x"f6",x"59",x"c6"),
   623 => (x"5b",x"5e",x"0e",x"87"),
   624 => (x"4a",x"71",x"0e",x"5c"),
   625 => (x"9a",x"72",x"4b",x"c0"),
   626 => (x"87",x"e1",x"c0",x"02"),
   627 => (x"9f",x"49",x"a2",x"da"),
   628 => (x"ea",x"c2",x"4b",x"69"),
   629 => (x"cf",x"02",x"bf",x"fe"),
   630 => (x"49",x"a2",x"d4",x"87"),
   631 => (x"4c",x"49",x"69",x"9f"),
   632 => (x"9c",x"ff",x"ff",x"c0"),
   633 => (x"87",x"c2",x"34",x"d0"),
   634 => (x"49",x"74",x"4c",x"c0"),
   635 => (x"fd",x"49",x"73",x"b3"),
   636 => (x"ef",x"f5",x"87",x"ed"),
   637 => (x"5b",x"5e",x"0e",x"87"),
   638 => (x"f4",x"0e",x"5d",x"5c"),
   639 => (x"c0",x"4a",x"71",x"86"),
   640 => (x"02",x"9a",x"72",x"7e"),
   641 => (x"e2",x"c2",x"87",x"d8"),
   642 => (x"78",x"c0",x"48",x"f2"),
   643 => (x"48",x"ea",x"e2",x"c2"),
   644 => (x"bf",x"e3",x"ef",x"c2"),
   645 => (x"ee",x"e2",x"c2",x"78"),
   646 => (x"df",x"ef",x"c2",x"48"),
   647 => (x"eb",x"c2",x"78",x"bf"),
   648 => (x"50",x"c0",x"48",x"d3"),
   649 => (x"bf",x"c2",x"eb",x"c2"),
   650 => (x"f2",x"e2",x"c2",x"49"),
   651 => (x"aa",x"71",x"4a",x"bf"),
   652 => (x"87",x"c9",x"c4",x"03"),
   653 => (x"99",x"cf",x"49",x"72"),
   654 => (x"87",x"e9",x"c0",x"05"),
   655 => (x"48",x"d0",x"ef",x"c0"),
   656 => (x"bf",x"ea",x"e2",x"c2"),
   657 => (x"f6",x"e2",x"c2",x"78"),
   658 => (x"ea",x"e2",x"c2",x"1e"),
   659 => (x"e2",x"c2",x"49",x"bf"),
   660 => (x"a1",x"c1",x"48",x"ea"),
   661 => (x"cb",x"e6",x"71",x"78"),
   662 => (x"c0",x"86",x"c4",x"87"),
   663 => (x"c2",x"48",x"cc",x"ef"),
   664 => (x"cc",x"78",x"f6",x"e2"),
   665 => (x"cc",x"ef",x"c0",x"87"),
   666 => (x"e0",x"c0",x"48",x"bf"),
   667 => (x"d0",x"ef",x"c0",x"80"),
   668 => (x"f2",x"e2",x"c2",x"58"),
   669 => (x"80",x"c1",x"48",x"bf"),
   670 => (x"58",x"f6",x"e2",x"c2"),
   671 => (x"00",x"0b",x"cc",x"27"),
   672 => (x"bf",x"97",x"bf",x"00"),
   673 => (x"c2",x"02",x"9d",x"4d"),
   674 => (x"e5",x"c3",x"87",x"e3"),
   675 => (x"dc",x"c2",x"02",x"ad"),
   676 => (x"cc",x"ef",x"c0",x"87"),
   677 => (x"a3",x"cb",x"4b",x"bf"),
   678 => (x"cf",x"4c",x"11",x"49"),
   679 => (x"d2",x"c1",x"05",x"ac"),
   680 => (x"df",x"49",x"75",x"87"),
   681 => (x"cd",x"89",x"c1",x"99"),
   682 => (x"c6",x"eb",x"c2",x"91"),
   683 => (x"4a",x"a3",x"c1",x"81"),
   684 => (x"a3",x"c3",x"51",x"12"),
   685 => (x"c5",x"51",x"12",x"4a"),
   686 => (x"51",x"12",x"4a",x"a3"),
   687 => (x"12",x"4a",x"a3",x"c7"),
   688 => (x"4a",x"a3",x"c9",x"51"),
   689 => (x"a3",x"ce",x"51",x"12"),
   690 => (x"d0",x"51",x"12",x"4a"),
   691 => (x"51",x"12",x"4a",x"a3"),
   692 => (x"12",x"4a",x"a3",x"d2"),
   693 => (x"4a",x"a3",x"d4",x"51"),
   694 => (x"a3",x"d6",x"51",x"12"),
   695 => (x"d8",x"51",x"12",x"4a"),
   696 => (x"51",x"12",x"4a",x"a3"),
   697 => (x"12",x"4a",x"a3",x"dc"),
   698 => (x"4a",x"a3",x"de",x"51"),
   699 => (x"7e",x"c1",x"51",x"12"),
   700 => (x"74",x"87",x"fa",x"c0"),
   701 => (x"05",x"99",x"c8",x"49"),
   702 => (x"74",x"87",x"eb",x"c0"),
   703 => (x"05",x"99",x"d0",x"49"),
   704 => (x"66",x"dc",x"87",x"d1"),
   705 => (x"87",x"cb",x"c0",x"02"),
   706 => (x"66",x"dc",x"49",x"73"),
   707 => (x"02",x"98",x"70",x"0f"),
   708 => (x"6e",x"87",x"d3",x"c0"),
   709 => (x"87",x"c6",x"c0",x"05"),
   710 => (x"48",x"c6",x"eb",x"c2"),
   711 => (x"ef",x"c0",x"50",x"c0"),
   712 => (x"c2",x"48",x"bf",x"cc"),
   713 => (x"eb",x"c2",x"87",x"e1"),
   714 => (x"50",x"c0",x"48",x"d3"),
   715 => (x"c2",x"eb",x"c2",x"7e"),
   716 => (x"e2",x"c2",x"49",x"bf"),
   717 => (x"71",x"4a",x"bf",x"f2"),
   718 => (x"f7",x"fb",x"04",x"aa"),
   719 => (x"e3",x"ef",x"c2",x"87"),
   720 => (x"c8",x"c0",x"05",x"bf"),
   721 => (x"fe",x"ea",x"c2",x"87"),
   722 => (x"f8",x"c1",x"02",x"bf"),
   723 => (x"ee",x"e2",x"c2",x"87"),
   724 => (x"d5",x"f0",x"49",x"bf"),
   725 => (x"c2",x"49",x"70",x"87"),
   726 => (x"c4",x"59",x"f2",x"e2"),
   727 => (x"e2",x"c2",x"48",x"a6"),
   728 => (x"c2",x"78",x"bf",x"ee"),
   729 => (x"02",x"bf",x"fe",x"ea"),
   730 => (x"c4",x"87",x"d8",x"c0"),
   731 => (x"ff",x"cf",x"49",x"66"),
   732 => (x"99",x"f8",x"ff",x"ff"),
   733 => (x"c5",x"c0",x"02",x"a9"),
   734 => (x"c0",x"4c",x"c0",x"87"),
   735 => (x"4c",x"c1",x"87",x"e1"),
   736 => (x"c4",x"87",x"dc",x"c0"),
   737 => (x"ff",x"cf",x"49",x"66"),
   738 => (x"02",x"a9",x"99",x"f8"),
   739 => (x"c8",x"87",x"c8",x"c0"),
   740 => (x"78",x"c0",x"48",x"a6"),
   741 => (x"c8",x"87",x"c5",x"c0"),
   742 => (x"78",x"c1",x"48",x"a6"),
   743 => (x"74",x"4c",x"66",x"c8"),
   744 => (x"e0",x"c0",x"05",x"9c"),
   745 => (x"49",x"66",x"c4",x"87"),
   746 => (x"ea",x"c2",x"89",x"c2"),
   747 => (x"91",x"4a",x"bf",x"f6"),
   748 => (x"bf",x"cf",x"ef",x"c2"),
   749 => (x"ea",x"e2",x"c2",x"4a"),
   750 => (x"78",x"a1",x"72",x"48"),
   751 => (x"48",x"f2",x"e2",x"c2"),
   752 => (x"df",x"f9",x"78",x"c0"),
   753 => (x"f4",x"48",x"c0",x"87"),
   754 => (x"87",x"d6",x"ee",x"8e"),
   755 => (x"00",x"00",x"00",x"00"),
   756 => (x"ff",x"ff",x"ff",x"ff"),
   757 => (x"00",x"00",x"0b",x"dc"),
   758 => (x"00",x"00",x"0b",x"e5"),
   759 => (x"33",x"54",x"41",x"46"),
   760 => (x"20",x"20",x"20",x"32"),
   761 => (x"54",x"41",x"46",x"00"),
   762 => (x"20",x"20",x"36",x"31"),
   763 => (x"ff",x"1e",x"00",x"20"),
   764 => (x"ff",x"c3",x"48",x"d4"),
   765 => (x"26",x"48",x"68",x"78"),
   766 => (x"d4",x"ff",x"1e",x"4f"),
   767 => (x"78",x"ff",x"c3",x"48"),
   768 => (x"c0",x"48",x"d0",x"ff"),
   769 => (x"d4",x"ff",x"78",x"e1"),
   770 => (x"c2",x"78",x"d4",x"48"),
   771 => (x"ff",x"48",x"e7",x"ef"),
   772 => (x"26",x"50",x"bf",x"d4"),
   773 => (x"d0",x"ff",x"1e",x"4f"),
   774 => (x"78",x"e0",x"c0",x"48"),
   775 => (x"ff",x"1e",x"4f",x"26"),
   776 => (x"49",x"70",x"87",x"cc"),
   777 => (x"87",x"c6",x"02",x"99"),
   778 => (x"05",x"a9",x"fb",x"c0"),
   779 => (x"48",x"71",x"87",x"f1"),
   780 => (x"5e",x"0e",x"4f",x"26"),
   781 => (x"71",x"0e",x"5c",x"5b"),
   782 => (x"fe",x"4c",x"c0",x"4b"),
   783 => (x"49",x"70",x"87",x"f0"),
   784 => (x"f9",x"c0",x"02",x"99"),
   785 => (x"a9",x"ec",x"c0",x"87"),
   786 => (x"87",x"f2",x"c0",x"02"),
   787 => (x"02",x"a9",x"fb",x"c0"),
   788 => (x"cc",x"87",x"eb",x"c0"),
   789 => (x"03",x"ac",x"b7",x"66"),
   790 => (x"66",x"d0",x"87",x"c7"),
   791 => (x"71",x"87",x"c2",x"02"),
   792 => (x"02",x"99",x"71",x"53"),
   793 => (x"84",x"c1",x"87",x"c2"),
   794 => (x"70",x"87",x"c3",x"fe"),
   795 => (x"cd",x"02",x"99",x"49"),
   796 => (x"a9",x"ec",x"c0",x"87"),
   797 => (x"c0",x"87",x"c7",x"02"),
   798 => (x"ff",x"05",x"a9",x"fb"),
   799 => (x"66",x"d0",x"87",x"d5"),
   800 => (x"c0",x"87",x"c3",x"02"),
   801 => (x"ec",x"c0",x"7b",x"97"),
   802 => (x"87",x"c4",x"05",x"a9"),
   803 => (x"87",x"c5",x"4a",x"74"),
   804 => (x"0a",x"c0",x"4a",x"74"),
   805 => (x"c2",x"48",x"72",x"8a"),
   806 => (x"26",x"4d",x"26",x"87"),
   807 => (x"26",x"4b",x"26",x"4c"),
   808 => (x"c9",x"fd",x"1e",x"4f"),
   809 => (x"4a",x"49",x"70",x"87"),
   810 => (x"04",x"aa",x"f0",x"c0"),
   811 => (x"f9",x"c0",x"87",x"c9"),
   812 => (x"87",x"c3",x"01",x"aa"),
   813 => (x"c1",x"8a",x"f0",x"c0"),
   814 => (x"c9",x"04",x"aa",x"c1"),
   815 => (x"aa",x"da",x"c1",x"87"),
   816 => (x"c0",x"87",x"c3",x"01"),
   817 => (x"48",x"72",x"8a",x"f7"),
   818 => (x"5e",x"0e",x"4f",x"26"),
   819 => (x"71",x"0e",x"5c",x"5b"),
   820 => (x"4b",x"d4",x"ff",x"4a"),
   821 => (x"e7",x"c0",x"49",x"72"),
   822 => (x"9c",x"4c",x"70",x"87"),
   823 => (x"c1",x"87",x"c2",x"02"),
   824 => (x"48",x"d0",x"ff",x"8c"),
   825 => (x"d5",x"c1",x"78",x"c5"),
   826 => (x"c6",x"49",x"74",x"7b"),
   827 => (x"c6",x"e0",x"c1",x"31"),
   828 => (x"48",x"4a",x"bf",x"97"),
   829 => (x"7b",x"70",x"b0",x"71"),
   830 => (x"c4",x"48",x"d0",x"ff"),
   831 => (x"87",x"db",x"fe",x"78"),
   832 => (x"5c",x"5b",x"5e",x"0e"),
   833 => (x"86",x"f8",x"0e",x"5d"),
   834 => (x"7e",x"c0",x"4c",x"71"),
   835 => (x"c0",x"87",x"ea",x"fb"),
   836 => (x"ed",x"f6",x"c0",x"4b"),
   837 => (x"c0",x"49",x"bf",x"97"),
   838 => (x"87",x"cf",x"04",x"a9"),
   839 => (x"c1",x"87",x"ff",x"fb"),
   840 => (x"ed",x"f6",x"c0",x"83"),
   841 => (x"ab",x"49",x"bf",x"97"),
   842 => (x"c0",x"87",x"f1",x"06"),
   843 => (x"bf",x"97",x"ed",x"f6"),
   844 => (x"fa",x"87",x"cf",x"02"),
   845 => (x"49",x"70",x"87",x"f8"),
   846 => (x"87",x"c6",x"02",x"99"),
   847 => (x"05",x"a9",x"ec",x"c0"),
   848 => (x"4b",x"c0",x"87",x"f1"),
   849 => (x"70",x"87",x"e7",x"fa"),
   850 => (x"87",x"e2",x"fa",x"4d"),
   851 => (x"fa",x"58",x"a6",x"c8"),
   852 => (x"4a",x"70",x"87",x"dc"),
   853 => (x"a4",x"c8",x"83",x"c1"),
   854 => (x"49",x"69",x"97",x"49"),
   855 => (x"87",x"c7",x"02",x"ad"),
   856 => (x"05",x"ad",x"ff",x"c0"),
   857 => (x"c9",x"87",x"e7",x"c0"),
   858 => (x"69",x"97",x"49",x"a4"),
   859 => (x"a9",x"66",x"c4",x"49"),
   860 => (x"48",x"87",x"c7",x"02"),
   861 => (x"05",x"a8",x"ff",x"c0"),
   862 => (x"a4",x"ca",x"87",x"d4"),
   863 => (x"49",x"69",x"97",x"49"),
   864 => (x"87",x"c6",x"02",x"aa"),
   865 => (x"05",x"aa",x"ff",x"c0"),
   866 => (x"7e",x"c1",x"87",x"c4"),
   867 => (x"ec",x"c0",x"87",x"d0"),
   868 => (x"87",x"c6",x"02",x"ad"),
   869 => (x"05",x"ad",x"fb",x"c0"),
   870 => (x"4b",x"c0",x"87",x"c4"),
   871 => (x"02",x"6e",x"7e",x"c1"),
   872 => (x"f9",x"87",x"e1",x"fe"),
   873 => (x"48",x"73",x"87",x"ef"),
   874 => (x"ec",x"fb",x"8e",x"f8"),
   875 => (x"5e",x"0e",x"00",x"87"),
   876 => (x"0e",x"5d",x"5c",x"5b"),
   877 => (x"4d",x"71",x"86",x"f8"),
   878 => (x"75",x"4b",x"d4",x"ff"),
   879 => (x"ec",x"ef",x"c2",x"1e"),
   880 => (x"87",x"d8",x"e8",x"49"),
   881 => (x"98",x"70",x"86",x"c4"),
   882 => (x"87",x"cc",x"c4",x"02"),
   883 => (x"c1",x"48",x"a6",x"c4"),
   884 => (x"78",x"bf",x"c8",x"e0"),
   885 => (x"f1",x"fb",x"49",x"75"),
   886 => (x"48",x"d0",x"ff",x"87"),
   887 => (x"d6",x"c1",x"78",x"c5"),
   888 => (x"75",x"4a",x"c0",x"7b"),
   889 => (x"7b",x"11",x"49",x"a2"),
   890 => (x"b7",x"cb",x"82",x"c1"),
   891 => (x"87",x"f3",x"04",x"aa"),
   892 => (x"ff",x"c3",x"4a",x"cc"),
   893 => (x"c0",x"82",x"c1",x"7b"),
   894 => (x"04",x"aa",x"b7",x"e0"),
   895 => (x"d0",x"ff",x"87",x"f4"),
   896 => (x"c3",x"78",x"c4",x"48"),
   897 => (x"78",x"c5",x"7b",x"ff"),
   898 => (x"c1",x"7b",x"d3",x"c1"),
   899 => (x"66",x"78",x"c4",x"7b"),
   900 => (x"a8",x"b7",x"c0",x"48"),
   901 => (x"87",x"f0",x"c2",x"06"),
   902 => (x"bf",x"f4",x"ef",x"c2"),
   903 => (x"48",x"66",x"c4",x"4c"),
   904 => (x"a6",x"c8",x"88",x"74"),
   905 => (x"02",x"9c",x"74",x"58"),
   906 => (x"c2",x"87",x"f9",x"c1"),
   907 => (x"c8",x"7e",x"f6",x"e2"),
   908 => (x"c0",x"8c",x"4d",x"c0"),
   909 => (x"c6",x"03",x"ac",x"b7"),
   910 => (x"a4",x"c0",x"c8",x"87"),
   911 => (x"c2",x"4c",x"c0",x"4d"),
   912 => (x"bf",x"97",x"e7",x"ef"),
   913 => (x"02",x"99",x"d0",x"49"),
   914 => (x"1e",x"c0",x"87",x"d1"),
   915 => (x"49",x"ec",x"ef",x"c2"),
   916 => (x"c4",x"87",x"fd",x"ea"),
   917 => (x"4a",x"49",x"70",x"86"),
   918 => (x"c2",x"87",x"ee",x"c0"),
   919 => (x"c2",x"1e",x"f6",x"e2"),
   920 => (x"ea",x"49",x"ec",x"ef"),
   921 => (x"86",x"c4",x"87",x"ea"),
   922 => (x"ff",x"4a",x"49",x"70"),
   923 => (x"c5",x"c8",x"48",x"d0"),
   924 => (x"7b",x"d4",x"c1",x"78"),
   925 => (x"7b",x"bf",x"97",x"6e"),
   926 => (x"80",x"c1",x"48",x"6e"),
   927 => (x"8d",x"c1",x"7e",x"70"),
   928 => (x"87",x"f0",x"ff",x"05"),
   929 => (x"c4",x"48",x"d0",x"ff"),
   930 => (x"05",x"9a",x"72",x"78"),
   931 => (x"48",x"c0",x"87",x"c5"),
   932 => (x"c1",x"87",x"c7",x"c1"),
   933 => (x"ec",x"ef",x"c2",x"1e"),
   934 => (x"87",x"da",x"e8",x"49"),
   935 => (x"9c",x"74",x"86",x"c4"),
   936 => (x"87",x"c7",x"fe",x"05"),
   937 => (x"c0",x"48",x"66",x"c4"),
   938 => (x"d1",x"06",x"a8",x"b7"),
   939 => (x"ec",x"ef",x"c2",x"87"),
   940 => (x"d0",x"78",x"c0",x"48"),
   941 => (x"f4",x"78",x"c0",x"80"),
   942 => (x"f8",x"ef",x"c2",x"80"),
   943 => (x"66",x"c4",x"78",x"bf"),
   944 => (x"a8",x"b7",x"c0",x"48"),
   945 => (x"87",x"d0",x"fd",x"01"),
   946 => (x"c5",x"48",x"d0",x"ff"),
   947 => (x"7b",x"d3",x"c1",x"78"),
   948 => (x"78",x"c4",x"7b",x"c0"),
   949 => (x"87",x"c2",x"48",x"c1"),
   950 => (x"8e",x"f8",x"48",x"c0"),
   951 => (x"4c",x"26",x"4d",x"26"),
   952 => (x"4f",x"26",x"4b",x"26"),
   953 => (x"5c",x"5b",x"5e",x"0e"),
   954 => (x"71",x"1e",x"0e",x"5d"),
   955 => (x"4d",x"4c",x"c0",x"4b"),
   956 => (x"e8",x"c0",x"04",x"ab"),
   957 => (x"c0",x"f4",x"c0",x"87"),
   958 => (x"02",x"9d",x"75",x"1e"),
   959 => (x"4a",x"c0",x"87",x"c4"),
   960 => (x"4a",x"c1",x"87",x"c2"),
   961 => (x"ec",x"eb",x"49",x"72"),
   962 => (x"70",x"86",x"c4",x"87"),
   963 => (x"6e",x"84",x"c1",x"7e"),
   964 => (x"73",x"87",x"c2",x"05"),
   965 => (x"73",x"85",x"c1",x"4c"),
   966 => (x"d8",x"ff",x"06",x"ac"),
   967 => (x"26",x"48",x"6e",x"87"),
   968 => (x"1e",x"87",x"f9",x"fe"),
   969 => (x"66",x"c4",x"4a",x"71"),
   970 => (x"72",x"87",x"c5",x"05"),
   971 => (x"87",x"fe",x"f9",x"49"),
   972 => (x"5e",x"0e",x"4f",x"26"),
   973 => (x"0e",x"5d",x"5c",x"5b"),
   974 => (x"49",x"4c",x"71",x"1e"),
   975 => (x"f0",x"c2",x"91",x"de"),
   976 => (x"85",x"71",x"4d",x"d4"),
   977 => (x"c1",x"02",x"6d",x"97"),
   978 => (x"f0",x"c2",x"87",x"dd"),
   979 => (x"74",x"4a",x"bf",x"c0"),
   980 => (x"fe",x"49",x"72",x"82"),
   981 => (x"7e",x"70",x"87",x"ce"),
   982 => (x"c0",x"02",x"98",x"48"),
   983 => (x"f0",x"c2",x"87",x"f2"),
   984 => (x"4a",x"70",x"4b",x"c8"),
   985 => (x"c4",x"ff",x"49",x"cb"),
   986 => (x"4b",x"74",x"87",x"fd"),
   987 => (x"e0",x"c1",x"93",x"cb"),
   988 => (x"83",x"c4",x"83",x"da"),
   989 => (x"7b",x"eb",x"fe",x"c0"),
   990 => (x"c1",x"c1",x"49",x"74"),
   991 => (x"7b",x"75",x"87",x"fd"),
   992 => (x"97",x"c7",x"e0",x"c1"),
   993 => (x"c2",x"1e",x"49",x"bf"),
   994 => (x"fe",x"49",x"c8",x"f0"),
   995 => (x"86",x"c4",x"87",x"d5"),
   996 => (x"c1",x"c1",x"49",x"74"),
   997 => (x"49",x"c0",x"87",x"e5"),
   998 => (x"87",x"c4",x"c3",x"c1"),
   999 => (x"48",x"e8",x"ef",x"c2"),
  1000 => (x"49",x"c1",x"78",x"c0"),
  1001 => (x"26",x"87",x"e6",x"dd"),
  1002 => (x"4c",x"87",x"f1",x"fc"),
  1003 => (x"69",x"64",x"61",x"6f"),
  1004 => (x"2e",x"2e",x"67",x"6e"),
  1005 => (x"5e",x"0e",x"00",x"2e"),
  1006 => (x"71",x"0e",x"5c",x"5b"),
  1007 => (x"f0",x"c2",x"4a",x"4b"),
  1008 => (x"72",x"82",x"bf",x"c0"),
  1009 => (x"87",x"dc",x"fc",x"49"),
  1010 => (x"02",x"9c",x"4c",x"70"),
  1011 => (x"e7",x"49",x"87",x"c4"),
  1012 => (x"f0",x"c2",x"87",x"eb"),
  1013 => (x"78",x"c0",x"48",x"c0"),
  1014 => (x"f0",x"dc",x"49",x"c1"),
  1015 => (x"87",x"fe",x"fb",x"87"),
  1016 => (x"5c",x"5b",x"5e",x"0e"),
  1017 => (x"86",x"f4",x"0e",x"5d"),
  1018 => (x"4d",x"f6",x"e2",x"c2"),
  1019 => (x"a6",x"c4",x"4c",x"c0"),
  1020 => (x"c2",x"78",x"c0",x"48"),
  1021 => (x"49",x"bf",x"c0",x"f0"),
  1022 => (x"c1",x"06",x"a9",x"c0"),
  1023 => (x"e2",x"c2",x"87",x"c1"),
  1024 => (x"02",x"98",x"48",x"f6"),
  1025 => (x"c0",x"87",x"f8",x"c0"),
  1026 => (x"c8",x"1e",x"c0",x"f4"),
  1027 => (x"87",x"c7",x"02",x"66"),
  1028 => (x"c0",x"48",x"a6",x"c4"),
  1029 => (x"c4",x"87",x"c5",x"78"),
  1030 => (x"78",x"c1",x"48",x"a6"),
  1031 => (x"e7",x"49",x"66",x"c4"),
  1032 => (x"86",x"c4",x"87",x"d3"),
  1033 => (x"84",x"c1",x"4d",x"70"),
  1034 => (x"c1",x"48",x"66",x"c4"),
  1035 => (x"58",x"a6",x"c8",x"80"),
  1036 => (x"bf",x"c0",x"f0",x"c2"),
  1037 => (x"c6",x"03",x"ac",x"49"),
  1038 => (x"05",x"9d",x"75",x"87"),
  1039 => (x"c0",x"87",x"c8",x"ff"),
  1040 => (x"02",x"9d",x"75",x"4c"),
  1041 => (x"c0",x"87",x"e0",x"c3"),
  1042 => (x"c8",x"1e",x"c0",x"f4"),
  1043 => (x"87",x"c7",x"02",x"66"),
  1044 => (x"c0",x"48",x"a6",x"cc"),
  1045 => (x"cc",x"87",x"c5",x"78"),
  1046 => (x"78",x"c1",x"48",x"a6"),
  1047 => (x"e6",x"49",x"66",x"cc"),
  1048 => (x"86",x"c4",x"87",x"d3"),
  1049 => (x"98",x"48",x"7e",x"70"),
  1050 => (x"87",x"e8",x"c2",x"02"),
  1051 => (x"97",x"81",x"cb",x"49"),
  1052 => (x"99",x"d0",x"49",x"69"),
  1053 => (x"87",x"d6",x"c1",x"02"),
  1054 => (x"4a",x"f6",x"fe",x"c0"),
  1055 => (x"91",x"cb",x"49",x"74"),
  1056 => (x"81",x"da",x"e0",x"c1"),
  1057 => (x"81",x"c8",x"79",x"72"),
  1058 => (x"74",x"51",x"ff",x"c3"),
  1059 => (x"c2",x"91",x"de",x"49"),
  1060 => (x"71",x"4d",x"d4",x"f0"),
  1061 => (x"97",x"c1",x"c2",x"85"),
  1062 => (x"49",x"a5",x"c1",x"7d"),
  1063 => (x"c2",x"51",x"e0",x"c0"),
  1064 => (x"bf",x"97",x"c6",x"eb"),
  1065 => (x"c1",x"87",x"d2",x"02"),
  1066 => (x"4b",x"a5",x"c2",x"84"),
  1067 => (x"4a",x"c6",x"eb",x"c2"),
  1068 => (x"ff",x"fe",x"49",x"db"),
  1069 => (x"db",x"c1",x"87",x"f1"),
  1070 => (x"49",x"a5",x"cd",x"87"),
  1071 => (x"84",x"c1",x"51",x"c0"),
  1072 => (x"6e",x"4b",x"a5",x"c2"),
  1073 => (x"fe",x"49",x"cb",x"4a"),
  1074 => (x"c1",x"87",x"dc",x"ff"),
  1075 => (x"fc",x"c0",x"87",x"c6"),
  1076 => (x"49",x"74",x"4a",x"f2"),
  1077 => (x"e0",x"c1",x"91",x"cb"),
  1078 => (x"79",x"72",x"81",x"da"),
  1079 => (x"97",x"c6",x"eb",x"c2"),
  1080 => (x"87",x"d8",x"02",x"bf"),
  1081 => (x"91",x"de",x"49",x"74"),
  1082 => (x"f0",x"c2",x"84",x"c1"),
  1083 => (x"83",x"71",x"4b",x"d4"),
  1084 => (x"4a",x"c6",x"eb",x"c2"),
  1085 => (x"fe",x"fe",x"49",x"dd"),
  1086 => (x"87",x"d8",x"87",x"ed"),
  1087 => (x"93",x"de",x"4b",x"74"),
  1088 => (x"83",x"d4",x"f0",x"c2"),
  1089 => (x"c0",x"49",x"a3",x"cb"),
  1090 => (x"73",x"84",x"c1",x"51"),
  1091 => (x"49",x"cb",x"4a",x"6e"),
  1092 => (x"87",x"d3",x"fe",x"fe"),
  1093 => (x"c1",x"48",x"66",x"c4"),
  1094 => (x"58",x"a6",x"c8",x"80"),
  1095 => (x"c0",x"03",x"ac",x"c7"),
  1096 => (x"05",x"6e",x"87",x"c5"),
  1097 => (x"74",x"87",x"e0",x"fc"),
  1098 => (x"f6",x"8e",x"f4",x"48"),
  1099 => (x"73",x"1e",x"87",x"ee"),
  1100 => (x"49",x"4b",x"71",x"1e"),
  1101 => (x"e0",x"c1",x"91",x"cb"),
  1102 => (x"a1",x"c8",x"81",x"da"),
  1103 => (x"c6",x"e0",x"c1",x"4a"),
  1104 => (x"c9",x"50",x"12",x"48"),
  1105 => (x"f6",x"c0",x"4a",x"a1"),
  1106 => (x"50",x"12",x"48",x"ed"),
  1107 => (x"e0",x"c1",x"81",x"ca"),
  1108 => (x"50",x"11",x"48",x"c7"),
  1109 => (x"97",x"c7",x"e0",x"c1"),
  1110 => (x"c0",x"1e",x"49",x"bf"),
  1111 => (x"87",x"c3",x"f7",x"49"),
  1112 => (x"48",x"e8",x"ef",x"c2"),
  1113 => (x"49",x"c1",x"78",x"de"),
  1114 => (x"26",x"87",x"e2",x"d6"),
  1115 => (x"1e",x"87",x"f1",x"f5"),
  1116 => (x"cb",x"49",x"4a",x"71"),
  1117 => (x"da",x"e0",x"c1",x"91"),
  1118 => (x"11",x"81",x"c8",x"81"),
  1119 => (x"ec",x"ef",x"c2",x"48"),
  1120 => (x"c0",x"f0",x"c2",x"58"),
  1121 => (x"c1",x"78",x"c0",x"48"),
  1122 => (x"87",x"c1",x"d6",x"49"),
  1123 => (x"c0",x"1e",x"4f",x"26"),
  1124 => (x"cb",x"fb",x"c0",x"49"),
  1125 => (x"1e",x"4f",x"26",x"87"),
  1126 => (x"d2",x"02",x"99",x"71"),
  1127 => (x"ef",x"e1",x"c1",x"87"),
  1128 => (x"f7",x"50",x"c0",x"48"),
  1129 => (x"ef",x"c5",x"c1",x"80"),
  1130 => (x"d3",x"e0",x"c1",x"40"),
  1131 => (x"c1",x"87",x"ce",x"78"),
  1132 => (x"c1",x"48",x"eb",x"e1"),
  1133 => (x"fc",x"78",x"cc",x"e0"),
  1134 => (x"ce",x"c6",x"c1",x"80"),
  1135 => (x"0e",x"4f",x"26",x"78"),
  1136 => (x"0e",x"5c",x"5b",x"5e"),
  1137 => (x"cb",x"4a",x"4c",x"71"),
  1138 => (x"da",x"e0",x"c1",x"92"),
  1139 => (x"49",x"a2",x"c8",x"82"),
  1140 => (x"97",x"4b",x"a2",x"c9"),
  1141 => (x"97",x"1e",x"4b",x"6b"),
  1142 => (x"ca",x"1e",x"49",x"69"),
  1143 => (x"c0",x"49",x"12",x"82"),
  1144 => (x"c0",x"87",x"c6",x"e6"),
  1145 => (x"87",x"e5",x"d4",x"49"),
  1146 => (x"f8",x"c0",x"49",x"74"),
  1147 => (x"8e",x"f8",x"87",x"cd"),
  1148 => (x"1e",x"87",x"eb",x"f3"),
  1149 => (x"4b",x"71",x"1e",x"73"),
  1150 => (x"87",x"c3",x"ff",x"49"),
  1151 => (x"fe",x"fe",x"49",x"73"),
  1152 => (x"c0",x"49",x"c0",x"87"),
  1153 => (x"f3",x"87",x"d9",x"f9"),
  1154 => (x"73",x"1e",x"87",x"d6"),
  1155 => (x"c6",x"4b",x"71",x"1e"),
  1156 => (x"db",x"02",x"4a",x"a3"),
  1157 => (x"02",x"8a",x"c1",x"87"),
  1158 => (x"02",x"8a",x"87",x"d6"),
  1159 => (x"8a",x"87",x"da",x"c1"),
  1160 => (x"87",x"fc",x"c0",x"02"),
  1161 => (x"e1",x"c0",x"02",x"8a"),
  1162 => (x"cb",x"02",x"8a",x"87"),
  1163 => (x"87",x"db",x"c1",x"87"),
  1164 => (x"fa",x"fc",x"49",x"c7"),
  1165 => (x"87",x"de",x"c1",x"87"),
  1166 => (x"bf",x"c0",x"f0",x"c2"),
  1167 => (x"87",x"cb",x"c1",x"02"),
  1168 => (x"c2",x"88",x"c1",x"48"),
  1169 => (x"c1",x"58",x"c4",x"f0"),
  1170 => (x"f0",x"c2",x"87",x"c1"),
  1171 => (x"c0",x"02",x"bf",x"c4"),
  1172 => (x"f0",x"c2",x"87",x"f9"),
  1173 => (x"c1",x"48",x"bf",x"c0"),
  1174 => (x"c4",x"f0",x"c2",x"80"),
  1175 => (x"87",x"eb",x"c0",x"58"),
  1176 => (x"bf",x"c0",x"f0",x"c2"),
  1177 => (x"c2",x"89",x"c6",x"49"),
  1178 => (x"c0",x"59",x"c4",x"f0"),
  1179 => (x"da",x"03",x"a9",x"b7"),
  1180 => (x"c0",x"f0",x"c2",x"87"),
  1181 => (x"d2",x"78",x"c0",x"48"),
  1182 => (x"c4",x"f0",x"c2",x"87"),
  1183 => (x"87",x"cb",x"02",x"bf"),
  1184 => (x"bf",x"c0",x"f0",x"c2"),
  1185 => (x"c2",x"80",x"c6",x"48"),
  1186 => (x"c0",x"58",x"c4",x"f0"),
  1187 => (x"87",x"fd",x"d1",x"49"),
  1188 => (x"f5",x"c0",x"49",x"73"),
  1189 => (x"c7",x"f1",x"87",x"e5"),
  1190 => (x"5b",x"5e",x"0e",x"87"),
  1191 => (x"ff",x"0e",x"5d",x"5c"),
  1192 => (x"a6",x"dc",x"86",x"d0"),
  1193 => (x"48",x"a6",x"c8",x"59"),
  1194 => (x"80",x"c4",x"78",x"c0"),
  1195 => (x"78",x"66",x"c4",x"c1"),
  1196 => (x"78",x"c1",x"80",x"c4"),
  1197 => (x"78",x"c1",x"80",x"c4"),
  1198 => (x"48",x"c4",x"f0",x"c2"),
  1199 => (x"ef",x"c2",x"78",x"c1"),
  1200 => (x"de",x"48",x"bf",x"e8"),
  1201 => (x"87",x"cb",x"05",x"a8"),
  1202 => (x"70",x"87",x"d5",x"f4"),
  1203 => (x"59",x"a6",x"cc",x"49"),
  1204 => (x"e4",x"87",x"f9",x"cf"),
  1205 => (x"c5",x"e5",x"87",x"e3"),
  1206 => (x"87",x"d2",x"e4",x"87"),
  1207 => (x"fb",x"c0",x"4c",x"70"),
  1208 => (x"fb",x"c1",x"02",x"ac"),
  1209 => (x"05",x"66",x"d8",x"87"),
  1210 => (x"c1",x"87",x"ed",x"c1"),
  1211 => (x"c4",x"4a",x"66",x"c0"),
  1212 => (x"72",x"7e",x"6a",x"82"),
  1213 => (x"c1",x"dc",x"c1",x"1e"),
  1214 => (x"49",x"66",x"c4",x"48"),
  1215 => (x"20",x"4a",x"a1",x"c8"),
  1216 => (x"05",x"aa",x"71",x"41"),
  1217 => (x"51",x"10",x"87",x"f9"),
  1218 => (x"c0",x"c1",x"4a",x"26"),
  1219 => (x"c4",x"c1",x"48",x"66"),
  1220 => (x"49",x"6a",x"78",x"ee"),
  1221 => (x"51",x"74",x"81",x"c7"),
  1222 => (x"49",x"66",x"c0",x"c1"),
  1223 => (x"51",x"c1",x"81",x"c8"),
  1224 => (x"49",x"66",x"c0",x"c1"),
  1225 => (x"51",x"c0",x"81",x"c9"),
  1226 => (x"49",x"66",x"c0",x"c1"),
  1227 => (x"51",x"c0",x"81",x"ca"),
  1228 => (x"1e",x"d8",x"1e",x"c1"),
  1229 => (x"81",x"c8",x"49",x"6a"),
  1230 => (x"c8",x"87",x"f7",x"e3"),
  1231 => (x"66",x"c4",x"c1",x"86"),
  1232 => (x"01",x"a8",x"c0",x"48"),
  1233 => (x"a6",x"c8",x"87",x"c7"),
  1234 => (x"ce",x"78",x"c1",x"48"),
  1235 => (x"66",x"c4",x"c1",x"87"),
  1236 => (x"d0",x"88",x"c1",x"48"),
  1237 => (x"87",x"c3",x"58",x"a6"),
  1238 => (x"d0",x"87",x"c3",x"e3"),
  1239 => (x"78",x"c2",x"48",x"a6"),
  1240 => (x"cd",x"02",x"9c",x"74"),
  1241 => (x"66",x"c8",x"87",x"e2"),
  1242 => (x"66",x"c8",x"c1",x"48"),
  1243 => (x"d7",x"cd",x"03",x"a8"),
  1244 => (x"48",x"a6",x"dc",x"87"),
  1245 => (x"80",x"e8",x"78",x"c0"),
  1246 => (x"f1",x"e1",x"78",x"c0"),
  1247 => (x"c1",x"4c",x"70",x"87"),
  1248 => (x"c2",x"05",x"ac",x"d0"),
  1249 => (x"66",x"c4",x"87",x"d7"),
  1250 => (x"87",x"d5",x"e4",x"7e"),
  1251 => (x"a6",x"c8",x"49",x"70"),
  1252 => (x"87",x"da",x"e1",x"59"),
  1253 => (x"ec",x"c0",x"4c",x"70"),
  1254 => (x"eb",x"c1",x"05",x"ac"),
  1255 => (x"49",x"66",x"c8",x"87"),
  1256 => (x"c0",x"c1",x"91",x"cb"),
  1257 => (x"a1",x"c4",x"81",x"66"),
  1258 => (x"c8",x"4d",x"6a",x"4a"),
  1259 => (x"66",x"c4",x"4a",x"a1"),
  1260 => (x"ef",x"c5",x"c1",x"52"),
  1261 => (x"87",x"f6",x"e0",x"79"),
  1262 => (x"02",x"9c",x"4c",x"70"),
  1263 => (x"fb",x"c0",x"87",x"d8"),
  1264 => (x"87",x"d2",x"02",x"ac"),
  1265 => (x"e5",x"e0",x"55",x"74"),
  1266 => (x"9c",x"4c",x"70",x"87"),
  1267 => (x"c0",x"87",x"c7",x"02"),
  1268 => (x"ff",x"05",x"ac",x"fb"),
  1269 => (x"e0",x"c0",x"87",x"ee"),
  1270 => (x"55",x"c1",x"c2",x"55"),
  1271 => (x"d8",x"7d",x"97",x"c0"),
  1272 => (x"a9",x"6e",x"49",x"66"),
  1273 => (x"c8",x"87",x"db",x"05"),
  1274 => (x"66",x"cc",x"48",x"66"),
  1275 => (x"87",x"ca",x"04",x"a8"),
  1276 => (x"c1",x"48",x"66",x"c8"),
  1277 => (x"58",x"a6",x"cc",x"80"),
  1278 => (x"66",x"cc",x"87",x"c8"),
  1279 => (x"d0",x"88",x"c1",x"48"),
  1280 => (x"df",x"ff",x"58",x"a6"),
  1281 => (x"4c",x"70",x"87",x"e8"),
  1282 => (x"05",x"ac",x"d0",x"c1"),
  1283 => (x"66",x"d4",x"87",x"c8"),
  1284 => (x"d8",x"80",x"c1",x"48"),
  1285 => (x"d0",x"c1",x"58",x"a6"),
  1286 => (x"e9",x"fd",x"02",x"ac"),
  1287 => (x"a6",x"e0",x"c0",x"87"),
  1288 => (x"78",x"66",x"d8",x"48"),
  1289 => (x"c0",x"48",x"66",x"c4"),
  1290 => (x"05",x"a8",x"66",x"e0"),
  1291 => (x"c0",x"87",x"eb",x"c9"),
  1292 => (x"c0",x"48",x"a6",x"e4"),
  1293 => (x"c0",x"48",x"74",x"78"),
  1294 => (x"7e",x"70",x"88",x"fb"),
  1295 => (x"c9",x"02",x"98",x"48"),
  1296 => (x"cb",x"48",x"87",x"ed"),
  1297 => (x"48",x"7e",x"70",x"88"),
  1298 => (x"cd",x"c1",x"02",x"98"),
  1299 => (x"88",x"c9",x"48",x"87"),
  1300 => (x"98",x"48",x"7e",x"70"),
  1301 => (x"87",x"c1",x"c4",x"02"),
  1302 => (x"70",x"88",x"c4",x"48"),
  1303 => (x"02",x"98",x"48",x"7e"),
  1304 => (x"c1",x"48",x"87",x"ce"),
  1305 => (x"48",x"7e",x"70",x"88"),
  1306 => (x"ec",x"c3",x"02",x"98"),
  1307 => (x"87",x"e1",x"c8",x"87"),
  1308 => (x"c0",x"48",x"a6",x"dc"),
  1309 => (x"dd",x"ff",x"78",x"f0"),
  1310 => (x"4c",x"70",x"87",x"f4"),
  1311 => (x"02",x"ac",x"ec",x"c0"),
  1312 => (x"c0",x"87",x"c4",x"c0"),
  1313 => (x"c0",x"5c",x"a6",x"e0"),
  1314 => (x"cd",x"02",x"ac",x"ec"),
  1315 => (x"dd",x"dd",x"ff",x"87"),
  1316 => (x"c0",x"4c",x"70",x"87"),
  1317 => (x"ff",x"05",x"ac",x"ec"),
  1318 => (x"ec",x"c0",x"87",x"f3"),
  1319 => (x"c4",x"c0",x"02",x"ac"),
  1320 => (x"c9",x"dd",x"ff",x"87"),
  1321 => (x"ca",x"1e",x"c0",x"87"),
  1322 => (x"49",x"66",x"d0",x"1e"),
  1323 => (x"c8",x"c1",x"91",x"cb"),
  1324 => (x"80",x"71",x"48",x"66"),
  1325 => (x"c8",x"58",x"a6",x"cc"),
  1326 => (x"80",x"c4",x"48",x"66"),
  1327 => (x"cc",x"58",x"a6",x"d0"),
  1328 => (x"ff",x"49",x"bf",x"66"),
  1329 => (x"c1",x"87",x"eb",x"dd"),
  1330 => (x"d4",x"1e",x"de",x"1e"),
  1331 => (x"ff",x"49",x"bf",x"66"),
  1332 => (x"d0",x"87",x"df",x"dd"),
  1333 => (x"c0",x"49",x"70",x"86"),
  1334 => (x"ec",x"c0",x"89",x"09"),
  1335 => (x"e8",x"c0",x"59",x"a6"),
  1336 => (x"a8",x"c0",x"48",x"66"),
  1337 => (x"87",x"ee",x"c0",x"06"),
  1338 => (x"48",x"66",x"e8",x"c0"),
  1339 => (x"c0",x"03",x"a8",x"dd"),
  1340 => (x"66",x"c4",x"87",x"e4"),
  1341 => (x"e8",x"c0",x"49",x"bf"),
  1342 => (x"e0",x"c0",x"81",x"66"),
  1343 => (x"66",x"e8",x"c0",x"51"),
  1344 => (x"c4",x"81",x"c1",x"49"),
  1345 => (x"c2",x"81",x"bf",x"66"),
  1346 => (x"e8",x"c0",x"51",x"c1"),
  1347 => (x"81",x"c2",x"49",x"66"),
  1348 => (x"81",x"bf",x"66",x"c4"),
  1349 => (x"48",x"6e",x"51",x"c0"),
  1350 => (x"78",x"ee",x"c4",x"c1"),
  1351 => (x"81",x"c8",x"49",x"6e"),
  1352 => (x"6e",x"51",x"66",x"d0"),
  1353 => (x"d4",x"81",x"c9",x"49"),
  1354 => (x"49",x"6e",x"51",x"66"),
  1355 => (x"66",x"dc",x"81",x"ca"),
  1356 => (x"48",x"66",x"d0",x"51"),
  1357 => (x"a6",x"d4",x"80",x"c1"),
  1358 => (x"48",x"66",x"c8",x"58"),
  1359 => (x"04",x"a8",x"66",x"cc"),
  1360 => (x"c8",x"87",x"cb",x"c0"),
  1361 => (x"80",x"c1",x"48",x"66"),
  1362 => (x"c5",x"58",x"a6",x"cc"),
  1363 => (x"66",x"cc",x"87",x"e1"),
  1364 => (x"d0",x"88",x"c1",x"48"),
  1365 => (x"d6",x"c5",x"58",x"a6"),
  1366 => (x"c4",x"dd",x"ff",x"87"),
  1367 => (x"c0",x"49",x"70",x"87"),
  1368 => (x"ff",x"59",x"a6",x"ec"),
  1369 => (x"70",x"87",x"fa",x"dc"),
  1370 => (x"a6",x"e0",x"c0",x"49"),
  1371 => (x"48",x"66",x"dc",x"59"),
  1372 => (x"05",x"a8",x"ec",x"c0"),
  1373 => (x"dc",x"87",x"ca",x"c0"),
  1374 => (x"e8",x"c0",x"48",x"a6"),
  1375 => (x"c4",x"c0",x"78",x"66"),
  1376 => (x"e9",x"d9",x"ff",x"87"),
  1377 => (x"49",x"66",x"c8",x"87"),
  1378 => (x"c0",x"c1",x"91",x"cb"),
  1379 => (x"80",x"71",x"48",x"66"),
  1380 => (x"c8",x"4a",x"7e",x"70"),
  1381 => (x"ca",x"49",x"6e",x"82"),
  1382 => (x"66",x"e8",x"c0",x"81"),
  1383 => (x"49",x"66",x"dc",x"51"),
  1384 => (x"e8",x"c0",x"81",x"c1"),
  1385 => (x"48",x"c1",x"89",x"66"),
  1386 => (x"49",x"70",x"30",x"71"),
  1387 => (x"97",x"71",x"89",x"c1"),
  1388 => (x"f0",x"f3",x"c2",x"7a"),
  1389 => (x"e8",x"c0",x"49",x"bf"),
  1390 => (x"6a",x"97",x"29",x"66"),
  1391 => (x"98",x"71",x"48",x"4a"),
  1392 => (x"58",x"a6",x"f0",x"c0"),
  1393 => (x"81",x"c4",x"49",x"6e"),
  1394 => (x"e0",x"c0",x"4d",x"69"),
  1395 => (x"66",x"c4",x"48",x"66"),
  1396 => (x"c8",x"c0",x"02",x"a8"),
  1397 => (x"48",x"a6",x"c4",x"87"),
  1398 => (x"c5",x"c0",x"78",x"c0"),
  1399 => (x"48",x"a6",x"c4",x"87"),
  1400 => (x"66",x"c4",x"78",x"c1"),
  1401 => (x"1e",x"e0",x"c0",x"1e"),
  1402 => (x"d9",x"ff",x"49",x"75"),
  1403 => (x"86",x"c8",x"87",x"c4"),
  1404 => (x"b7",x"c0",x"4c",x"70"),
  1405 => (x"d4",x"c1",x"06",x"ac"),
  1406 => (x"c0",x"85",x"74",x"87"),
  1407 => (x"89",x"74",x"49",x"e0"),
  1408 => (x"dc",x"c1",x"4b",x"75"),
  1409 => (x"fe",x"71",x"4a",x"ca"),
  1410 => (x"c2",x"87",x"dc",x"ea"),
  1411 => (x"66",x"e4",x"c0",x"85"),
  1412 => (x"c0",x"80",x"c1",x"48"),
  1413 => (x"c0",x"58",x"a6",x"e8"),
  1414 => (x"c1",x"49",x"66",x"ec"),
  1415 => (x"02",x"a9",x"70",x"81"),
  1416 => (x"c4",x"87",x"c8",x"c0"),
  1417 => (x"78",x"c0",x"48",x"a6"),
  1418 => (x"c4",x"87",x"c5",x"c0"),
  1419 => (x"78",x"c1",x"48",x"a6"),
  1420 => (x"c2",x"1e",x"66",x"c4"),
  1421 => (x"e0",x"c0",x"49",x"a4"),
  1422 => (x"70",x"88",x"71",x"48"),
  1423 => (x"49",x"75",x"1e",x"49"),
  1424 => (x"87",x"ee",x"d7",x"ff"),
  1425 => (x"b7",x"c0",x"86",x"c8"),
  1426 => (x"c0",x"ff",x"01",x"a8"),
  1427 => (x"66",x"e4",x"c0",x"87"),
  1428 => (x"87",x"d1",x"c0",x"02"),
  1429 => (x"81",x"c9",x"49",x"6e"),
  1430 => (x"51",x"66",x"e4",x"c0"),
  1431 => (x"c6",x"c1",x"48",x"6e"),
  1432 => (x"cc",x"c0",x"78",x"ff"),
  1433 => (x"c9",x"49",x"6e",x"87"),
  1434 => (x"6e",x"51",x"c2",x"81"),
  1435 => (x"f3",x"c7",x"c1",x"48"),
  1436 => (x"48",x"66",x"c8",x"78"),
  1437 => (x"04",x"a8",x"66",x"cc"),
  1438 => (x"c8",x"87",x"cb",x"c0"),
  1439 => (x"80",x"c1",x"48",x"66"),
  1440 => (x"c0",x"58",x"a6",x"cc"),
  1441 => (x"66",x"cc",x"87",x"e9"),
  1442 => (x"d0",x"88",x"c1",x"48"),
  1443 => (x"de",x"c0",x"58",x"a6"),
  1444 => (x"c9",x"d6",x"ff",x"87"),
  1445 => (x"c0",x"4c",x"70",x"87"),
  1446 => (x"c6",x"c1",x"87",x"d5"),
  1447 => (x"c8",x"c0",x"05",x"ac"),
  1448 => (x"48",x"66",x"d0",x"87"),
  1449 => (x"a6",x"d4",x"80",x"c1"),
  1450 => (x"f1",x"d5",x"ff",x"58"),
  1451 => (x"d4",x"4c",x"70",x"87"),
  1452 => (x"80",x"c1",x"48",x"66"),
  1453 => (x"74",x"58",x"a6",x"d8"),
  1454 => (x"cb",x"c0",x"02",x"9c"),
  1455 => (x"48",x"66",x"c8",x"87"),
  1456 => (x"a8",x"66",x"c8",x"c1"),
  1457 => (x"87",x"e9",x"f2",x"04"),
  1458 => (x"87",x"c9",x"d5",x"ff"),
  1459 => (x"c7",x"48",x"66",x"c8"),
  1460 => (x"e5",x"c0",x"03",x"a8"),
  1461 => (x"c4",x"f0",x"c2",x"87"),
  1462 => (x"c8",x"78",x"c0",x"48"),
  1463 => (x"91",x"cb",x"49",x"66"),
  1464 => (x"81",x"66",x"c0",x"c1"),
  1465 => (x"6a",x"4a",x"a1",x"c4"),
  1466 => (x"79",x"52",x"c0",x"4a"),
  1467 => (x"c1",x"48",x"66",x"c8"),
  1468 => (x"58",x"a6",x"cc",x"80"),
  1469 => (x"ff",x"04",x"a8",x"c7"),
  1470 => (x"d0",x"ff",x"87",x"db"),
  1471 => (x"db",x"df",x"ff",x"8e"),
  1472 => (x"61",x"6f",x"4c",x"87"),
  1473 => (x"2e",x"2a",x"20",x"64"),
  1474 => (x"20",x"3a",x"00",x"20"),
  1475 => (x"1e",x"73",x"1e",x"00"),
  1476 => (x"02",x"9b",x"4b",x"71"),
  1477 => (x"f0",x"c2",x"87",x"c6"),
  1478 => (x"78",x"c0",x"48",x"c0"),
  1479 => (x"f0",x"c2",x"1e",x"c7"),
  1480 => (x"1e",x"49",x"bf",x"c0"),
  1481 => (x"1e",x"da",x"e0",x"c1"),
  1482 => (x"bf",x"e8",x"ef",x"c2"),
  1483 => (x"87",x"e9",x"ed",x"49"),
  1484 => (x"ef",x"c2",x"86",x"cc"),
  1485 => (x"e9",x"49",x"bf",x"e8"),
  1486 => (x"9b",x"73",x"87",x"dd"),
  1487 => (x"c1",x"87",x"c8",x"02"),
  1488 => (x"c0",x"49",x"da",x"e0"),
  1489 => (x"ff",x"87",x"c6",x"e4"),
  1490 => (x"1e",x"87",x"d5",x"de"),
  1491 => (x"4b",x"c0",x"1e",x"73"),
  1492 => (x"48",x"c6",x"e0",x"c1"),
  1493 => (x"e1",x"c1",x"50",x"c0"),
  1494 => (x"ff",x"49",x"bf",x"fd"),
  1495 => (x"70",x"87",x"cf",x"d9"),
  1496 => (x"87",x"c4",x"05",x"98"),
  1497 => (x"4b",x"ee",x"dd",x"c1"),
  1498 => (x"dd",x"ff",x"48",x"73"),
  1499 => (x"4f",x"52",x"87",x"f2"),
  1500 => (x"6f",x"6c",x"20",x"4d"),
  1501 => (x"6e",x"69",x"64",x"61"),
  1502 => (x"61",x"66",x"20",x"67"),
  1503 => (x"64",x"65",x"6c",x"69"),
  1504 => (x"df",x"c7",x"1e",x"00"),
  1505 => (x"fe",x"49",x"c1",x"87"),
  1506 => (x"ed",x"fe",x"87",x"c3"),
  1507 => (x"98",x"70",x"87",x"ff"),
  1508 => (x"fe",x"87",x"cd",x"02"),
  1509 => (x"70",x"87",x"d8",x"f5"),
  1510 => (x"87",x"c4",x"02",x"98"),
  1511 => (x"87",x"c2",x"4a",x"c1"),
  1512 => (x"9a",x"72",x"4a",x"c0"),
  1513 => (x"c0",x"87",x"ce",x"05"),
  1514 => (x"d1",x"df",x"c1",x"1e"),
  1515 => (x"d4",x"ef",x"c0",x"49"),
  1516 => (x"fe",x"86",x"c4",x"87"),
  1517 => (x"c1",x"1e",x"c0",x"87"),
  1518 => (x"c0",x"49",x"dc",x"df"),
  1519 => (x"c0",x"87",x"c6",x"ef"),
  1520 => (x"87",x"c7",x"fe",x"1e"),
  1521 => (x"ee",x"c0",x"49",x"70"),
  1522 => (x"d6",x"c3",x"87",x"fb"),
  1523 => (x"26",x"8e",x"f8",x"87"),
  1524 => (x"20",x"44",x"53",x"4f"),
  1525 => (x"6c",x"69",x"61",x"66"),
  1526 => (x"00",x"2e",x"64",x"65"),
  1527 => (x"74",x"6f",x"6f",x"42"),
  1528 => (x"2e",x"67",x"6e",x"69"),
  1529 => (x"1e",x"00",x"2e",x"2e"),
  1530 => (x"87",x"df",x"e6",x"c0"),
  1531 => (x"4f",x"26",x"87",x"fa"),
  1532 => (x"c0",x"f0",x"c2",x"1e"),
  1533 => (x"c2",x"78",x"c0",x"48"),
  1534 => (x"c0",x"48",x"e8",x"ef"),
  1535 => (x"87",x"c1",x"fe",x"78"),
  1536 => (x"48",x"c0",x"87",x"e5"),
  1537 => (x"00",x"00",x"4f",x"26"),
  1538 => (x"00",x"00",x"00",x"01"),
  1539 => (x"78",x"45",x"20",x"80"),
  1540 => (x"80",x"00",x"74",x"69"),
  1541 => (x"63",x"61",x"42",x"20"),
  1542 => (x"0f",x"32",x"00",x"6b"),
  1543 => (x"2c",x"14",x"00",x"00"),
  1544 => (x"00",x"00",x"00",x"00"),
  1545 => (x"00",x"0f",x"32",x"00"),
  1546 => (x"00",x"2c",x"32",x"00"),
  1547 => (x"00",x"00",x"00",x"00"),
  1548 => (x"00",x"00",x"0f",x"32"),
  1549 => (x"00",x"00",x"2c",x"50"),
  1550 => (x"32",x"00",x"00",x"00"),
  1551 => (x"6e",x"00",x"00",x"0f"),
  1552 => (x"00",x"00",x"00",x"2c"),
  1553 => (x"0f",x"32",x"00",x"00"),
  1554 => (x"2c",x"8c",x"00",x"00"),
  1555 => (x"00",x"00",x"00",x"00"),
  1556 => (x"00",x"0f",x"32",x"00"),
  1557 => (x"00",x"2c",x"aa",x"00"),
  1558 => (x"00",x"00",x"00",x"00"),
  1559 => (x"00",x"00",x"0f",x"32"),
  1560 => (x"00",x"00",x"2c",x"c8"),
  1561 => (x"6f",x"00",x"00",x"00"),
  1562 => (x"00",x"00",x"00",x"11"),
  1563 => (x"00",x"00",x"00",x"00"),
  1564 => (x"12",x"0a",x"00",x"00"),
  1565 => (x"00",x"00",x"00",x"00"),
  1566 => (x"00",x"00",x"00",x"00"),
  1567 => (x"00",x"18",x"81",x"00"),
  1568 => (x"54",x"45",x"50",x"00"),
  1569 => (x"31",x"30",x"30",x"32"),
  1570 => (x"4d",x"4f",x"52",x"20"),
  1571 => (x"f0",x"fe",x"1e",x"00"),
  1572 => (x"cd",x"78",x"c0",x"48"),
  1573 => (x"26",x"09",x"79",x"09"),
  1574 => (x"fe",x"1e",x"1e",x"4f"),
  1575 => (x"48",x"7e",x"bf",x"f0"),
  1576 => (x"1e",x"4f",x"26",x"26"),
  1577 => (x"c1",x"48",x"f0",x"fe"),
  1578 => (x"1e",x"4f",x"26",x"78"),
  1579 => (x"c0",x"48",x"f0",x"fe"),
  1580 => (x"1e",x"4f",x"26",x"78"),
  1581 => (x"52",x"c0",x"4a",x"71"),
  1582 => (x"0e",x"4f",x"26",x"52"),
  1583 => (x"5d",x"5c",x"5b",x"5e"),
  1584 => (x"71",x"86",x"f4",x"0e"),
  1585 => (x"7e",x"6d",x"97",x"4d"),
  1586 => (x"97",x"4c",x"a5",x"c1"),
  1587 => (x"a6",x"c8",x"48",x"6c"),
  1588 => (x"c4",x"48",x"6e",x"58"),
  1589 => (x"c5",x"05",x"a8",x"66"),
  1590 => (x"c0",x"48",x"ff",x"87"),
  1591 => (x"ca",x"ff",x"87",x"e6"),
  1592 => (x"49",x"a5",x"c2",x"87"),
  1593 => (x"71",x"4b",x"6c",x"97"),
  1594 => (x"6b",x"97",x"4b",x"a3"),
  1595 => (x"7e",x"6c",x"97",x"4b"),
  1596 => (x"80",x"c1",x"48",x"6e"),
  1597 => (x"c7",x"58",x"a6",x"c8"),
  1598 => (x"58",x"a6",x"cc",x"98"),
  1599 => (x"fe",x"7c",x"97",x"70"),
  1600 => (x"48",x"73",x"87",x"e1"),
  1601 => (x"4d",x"26",x"8e",x"f4"),
  1602 => (x"4b",x"26",x"4c",x"26"),
  1603 => (x"5e",x"0e",x"4f",x"26"),
  1604 => (x"f4",x"0e",x"5c",x"5b"),
  1605 => (x"d8",x"4c",x"71",x"86"),
  1606 => (x"ff",x"c3",x"4a",x"66"),
  1607 => (x"4b",x"a4",x"c2",x"9a"),
  1608 => (x"73",x"49",x"6c",x"97"),
  1609 => (x"51",x"72",x"49",x"a1"),
  1610 => (x"6e",x"7e",x"6c",x"97"),
  1611 => (x"c8",x"80",x"c1",x"48"),
  1612 => (x"98",x"c7",x"58",x"a6"),
  1613 => (x"70",x"58",x"a6",x"cc"),
  1614 => (x"ff",x"8e",x"f4",x"54"),
  1615 => (x"1e",x"1e",x"87",x"ca"),
  1616 => (x"e0",x"87",x"e8",x"fd"),
  1617 => (x"c0",x"49",x"4a",x"bf"),
  1618 => (x"02",x"99",x"c0",x"e0"),
  1619 => (x"1e",x"72",x"87",x"cb"),
  1620 => (x"49",x"e6",x"f3",x"c2"),
  1621 => (x"c4",x"87",x"f7",x"fe"),
  1622 => (x"87",x"fd",x"fc",x"86"),
  1623 => (x"c2",x"fd",x"7e",x"70"),
  1624 => (x"4f",x"26",x"26",x"87"),
  1625 => (x"e6",x"f3",x"c2",x"1e"),
  1626 => (x"87",x"c7",x"fd",x"49"),
  1627 => (x"49",x"fe",x"e4",x"c1"),
  1628 => (x"c3",x"87",x"da",x"fc"),
  1629 => (x"4f",x"26",x"87",x"ee"),
  1630 => (x"5c",x"5b",x"5e",x"0e"),
  1631 => (x"4d",x"71",x"0e",x"5d"),
  1632 => (x"49",x"e6",x"f3",x"c2"),
  1633 => (x"70",x"87",x"f4",x"fc"),
  1634 => (x"ab",x"b7",x"c0",x"4b"),
  1635 => (x"87",x"c2",x"c3",x"04"),
  1636 => (x"05",x"ab",x"f0",x"c3"),
  1637 => (x"e9",x"c1",x"87",x"c9"),
  1638 => (x"78",x"c1",x"48",x"dc"),
  1639 => (x"c3",x"87",x"e3",x"c2"),
  1640 => (x"c9",x"05",x"ab",x"e0"),
  1641 => (x"e0",x"e9",x"c1",x"87"),
  1642 => (x"c2",x"78",x"c1",x"48"),
  1643 => (x"e9",x"c1",x"87",x"d4"),
  1644 => (x"c6",x"02",x"bf",x"e0"),
  1645 => (x"a3",x"c0",x"c2",x"87"),
  1646 => (x"73",x"87",x"c2",x"4c"),
  1647 => (x"dc",x"e9",x"c1",x"4c"),
  1648 => (x"e0",x"c0",x"02",x"bf"),
  1649 => (x"c4",x"49",x"74",x"87"),
  1650 => (x"c1",x"91",x"29",x"b7"),
  1651 => (x"74",x"81",x"f3",x"ea"),
  1652 => (x"c2",x"9a",x"cf",x"4a"),
  1653 => (x"72",x"48",x"c1",x"92"),
  1654 => (x"ff",x"4a",x"70",x"30"),
  1655 => (x"69",x"48",x"72",x"ba"),
  1656 => (x"db",x"79",x"70",x"98"),
  1657 => (x"c4",x"49",x"74",x"87"),
  1658 => (x"c1",x"91",x"29",x"b7"),
  1659 => (x"74",x"81",x"f3",x"ea"),
  1660 => (x"c2",x"9a",x"cf",x"4a"),
  1661 => (x"72",x"48",x"c3",x"92"),
  1662 => (x"48",x"4a",x"70",x"30"),
  1663 => (x"79",x"70",x"b0",x"69"),
  1664 => (x"c0",x"05",x"9d",x"75"),
  1665 => (x"d0",x"ff",x"87",x"f0"),
  1666 => (x"78",x"e1",x"c8",x"48"),
  1667 => (x"c5",x"48",x"d4",x"ff"),
  1668 => (x"e0",x"e9",x"c1",x"78"),
  1669 => (x"87",x"c3",x"02",x"bf"),
  1670 => (x"c1",x"78",x"e0",x"c3"),
  1671 => (x"02",x"bf",x"dc",x"e9"),
  1672 => (x"d4",x"ff",x"87",x"c6"),
  1673 => (x"78",x"f0",x"c3",x"48"),
  1674 => (x"73",x"48",x"d4",x"ff"),
  1675 => (x"48",x"d0",x"ff",x"78"),
  1676 => (x"c0",x"78",x"e1",x"c8"),
  1677 => (x"e9",x"c1",x"78",x"e0"),
  1678 => (x"78",x"c0",x"48",x"e0"),
  1679 => (x"48",x"dc",x"e9",x"c1"),
  1680 => (x"f3",x"c2",x"78",x"c0"),
  1681 => (x"f2",x"f9",x"49",x"e6"),
  1682 => (x"c0",x"4b",x"70",x"87"),
  1683 => (x"fc",x"03",x"ab",x"b7"),
  1684 => (x"48",x"c0",x"87",x"fe"),
  1685 => (x"4c",x"26",x"4d",x"26"),
  1686 => (x"4f",x"26",x"4b",x"26"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"72",x"4a",x"c0",x"1e"),
  1690 => (x"c1",x"91",x"c4",x"49"),
  1691 => (x"c0",x"81",x"f3",x"ea"),
  1692 => (x"d0",x"82",x"c1",x"79"),
  1693 => (x"ee",x"04",x"aa",x"b7"),
  1694 => (x"0e",x"4f",x"26",x"87"),
  1695 => (x"5d",x"5c",x"5b",x"5e"),
  1696 => (x"f8",x"4d",x"71",x"0e"),
  1697 => (x"4a",x"75",x"87",x"e5"),
  1698 => (x"92",x"2a",x"b7",x"c4"),
  1699 => (x"82",x"f3",x"ea",x"c1"),
  1700 => (x"9c",x"cf",x"4c",x"75"),
  1701 => (x"49",x"6a",x"94",x"c2"),
  1702 => (x"c3",x"2b",x"74",x"4b"),
  1703 => (x"74",x"48",x"c2",x"9b"),
  1704 => (x"ff",x"4c",x"70",x"30"),
  1705 => (x"71",x"48",x"74",x"bc"),
  1706 => (x"f7",x"7a",x"70",x"98"),
  1707 => (x"48",x"73",x"87",x"f5"),
  1708 => (x"00",x"87",x"e1",x"fe"),
  1709 => (x"00",x"00",x"00",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"00",x"00"),
  1712 => (x"00",x"00",x"00",x"00"),
  1713 => (x"00",x"00",x"00",x"00"),
  1714 => (x"00",x"00",x"00",x"00"),
  1715 => (x"00",x"00",x"00",x"00"),
  1716 => (x"00",x"00",x"00",x"00"),
  1717 => (x"00",x"00",x"00",x"00"),
  1718 => (x"00",x"00",x"00",x"00"),
  1719 => (x"00",x"00",x"00",x"00"),
  1720 => (x"00",x"00",x"00",x"00"),
  1721 => (x"00",x"00",x"00",x"00"),
  1722 => (x"00",x"00",x"00",x"00"),
  1723 => (x"00",x"00",x"00",x"00"),
  1724 => (x"1e",x"00",x"00",x"00"),
  1725 => (x"c8",x"48",x"d0",x"ff"),
  1726 => (x"48",x"71",x"78",x"e1"),
  1727 => (x"78",x"08",x"d4",x"ff"),
  1728 => (x"ff",x"48",x"66",x"c4"),
  1729 => (x"26",x"78",x"08",x"d4"),
  1730 => (x"4a",x"71",x"1e",x"4f"),
  1731 => (x"1e",x"49",x"66",x"c4"),
  1732 => (x"de",x"ff",x"49",x"72"),
  1733 => (x"48",x"d0",x"ff",x"87"),
  1734 => (x"26",x"78",x"e0",x"c0"),
  1735 => (x"73",x"1e",x"4f",x"26"),
  1736 => (x"c8",x"4b",x"71",x"1e"),
  1737 => (x"73",x"1e",x"49",x"66"),
  1738 => (x"a2",x"e0",x"c1",x"4a"),
  1739 => (x"87",x"d9",x"ff",x"49"),
  1740 => (x"26",x"87",x"c4",x"26"),
  1741 => (x"26",x"4c",x"26",x"4d"),
  1742 => (x"1e",x"4f",x"26",x"4b"),
  1743 => (x"c3",x"4a",x"d4",x"ff"),
  1744 => (x"d0",x"ff",x"7a",x"ff"),
  1745 => (x"78",x"e1",x"c0",x"48"),
  1746 => (x"f3",x"c2",x"7a",x"de"),
  1747 => (x"49",x"7a",x"bf",x"f0"),
  1748 => (x"70",x"28",x"c8",x"48"),
  1749 => (x"d0",x"48",x"71",x"7a"),
  1750 => (x"71",x"7a",x"70",x"28"),
  1751 => (x"70",x"28",x"d8",x"48"),
  1752 => (x"48",x"d0",x"ff",x"7a"),
  1753 => (x"26",x"78",x"e0",x"c0"),
  1754 => (x"5b",x"5e",x"0e",x"4f"),
  1755 => (x"71",x"0e",x"5d",x"5c"),
  1756 => (x"f0",x"f3",x"c2",x"4c"),
  1757 => (x"74",x"49",x"4d",x"bf"),
  1758 => (x"d0",x"4b",x"71",x"29"),
  1759 => (x"83",x"c1",x"9b",x"66"),
  1760 => (x"ab",x"b7",x"66",x"d4"),
  1761 => (x"c0",x"87",x"c2",x"04"),
  1762 => (x"49",x"66",x"d0",x"4b"),
  1763 => (x"b9",x"ff",x"31",x"74"),
  1764 => (x"4a",x"73",x"99",x"75"),
  1765 => (x"48",x"72",x"32",x"74"),
  1766 => (x"f3",x"c2",x"b0",x"71"),
  1767 => (x"da",x"fe",x"58",x"f4"),
  1768 => (x"26",x"4d",x"26",x"87"),
  1769 => (x"26",x"4b",x"26",x"4c"),
  1770 => (x"d0",x"ff",x"1e",x"4f"),
  1771 => (x"78",x"c9",x"c8",x"48"),
  1772 => (x"d4",x"ff",x"48",x"71"),
  1773 => (x"4f",x"26",x"78",x"08"),
  1774 => (x"49",x"4a",x"71",x"1e"),
  1775 => (x"d0",x"ff",x"87",x"eb"),
  1776 => (x"26",x"78",x"c8",x"48"),
  1777 => (x"1e",x"73",x"1e",x"4f"),
  1778 => (x"f4",x"c2",x"4b",x"71"),
  1779 => (x"c3",x"02",x"bf",x"c0"),
  1780 => (x"87",x"eb",x"c2",x"87"),
  1781 => (x"c8",x"48",x"d0",x"ff"),
  1782 => (x"49",x"73",x"78",x"c9"),
  1783 => (x"ff",x"b1",x"e0",x"c0"),
  1784 => (x"78",x"71",x"48",x"d4"),
  1785 => (x"48",x"f4",x"f3",x"c2"),
  1786 => (x"66",x"c8",x"78",x"c0"),
  1787 => (x"c3",x"87",x"c5",x"02"),
  1788 => (x"87",x"c2",x"49",x"ff"),
  1789 => (x"f3",x"c2",x"49",x"c0"),
  1790 => (x"66",x"cc",x"59",x"fc"),
  1791 => (x"c5",x"87",x"c6",x"02"),
  1792 => (x"c4",x"4a",x"d5",x"d5"),
  1793 => (x"ff",x"ff",x"cf",x"87"),
  1794 => (x"c0",x"f4",x"c2",x"4a"),
  1795 => (x"c0",x"f4",x"c2",x"5a"),
  1796 => (x"c4",x"78",x"c1",x"48"),
  1797 => (x"26",x"4d",x"26",x"87"),
  1798 => (x"26",x"4b",x"26",x"4c"),
  1799 => (x"5b",x"5e",x"0e",x"4f"),
  1800 => (x"71",x"0e",x"5d",x"5c"),
  1801 => (x"fc",x"f3",x"c2",x"4a"),
  1802 => (x"9a",x"72",x"4c",x"bf"),
  1803 => (x"49",x"87",x"cb",x"02"),
  1804 => (x"ee",x"c1",x"91",x"c8"),
  1805 => (x"83",x"71",x"4b",x"fb"),
  1806 => (x"f2",x"c1",x"87",x"c4"),
  1807 => (x"4d",x"c0",x"4b",x"fb"),
  1808 => (x"99",x"74",x"49",x"13"),
  1809 => (x"bf",x"f8",x"f3",x"c2"),
  1810 => (x"48",x"d4",x"ff",x"b9"),
  1811 => (x"b7",x"c1",x"78",x"71"),
  1812 => (x"b7",x"c8",x"85",x"2c"),
  1813 => (x"87",x"e8",x"04",x"ad"),
  1814 => (x"bf",x"f4",x"f3",x"c2"),
  1815 => (x"c2",x"80",x"c8",x"48"),
  1816 => (x"fe",x"58",x"f8",x"f3"),
  1817 => (x"73",x"1e",x"87",x"ef"),
  1818 => (x"13",x"4b",x"71",x"1e"),
  1819 => (x"cb",x"02",x"9a",x"4a"),
  1820 => (x"fe",x"49",x"72",x"87"),
  1821 => (x"4a",x"13",x"87",x"e7"),
  1822 => (x"87",x"f5",x"05",x"9a"),
  1823 => (x"1e",x"87",x"da",x"fe"),
  1824 => (x"bf",x"f4",x"f3",x"c2"),
  1825 => (x"f4",x"f3",x"c2",x"49"),
  1826 => (x"78",x"a1",x"c1",x"48"),
  1827 => (x"a9",x"b7",x"c0",x"c4"),
  1828 => (x"ff",x"87",x"db",x"03"),
  1829 => (x"f3",x"c2",x"48",x"d4"),
  1830 => (x"c2",x"78",x"bf",x"f8"),
  1831 => (x"49",x"bf",x"f4",x"f3"),
  1832 => (x"48",x"f4",x"f3",x"c2"),
  1833 => (x"c4",x"78",x"a1",x"c1"),
  1834 => (x"04",x"a9",x"b7",x"c0"),
  1835 => (x"d0",x"ff",x"87",x"e5"),
  1836 => (x"c2",x"78",x"c8",x"48"),
  1837 => (x"c0",x"48",x"c0",x"f4"),
  1838 => (x"00",x"4f",x"26",x"78"),
  1839 => (x"00",x"00",x"00",x"00"),
  1840 => (x"00",x"00",x"00",x"00"),
  1841 => (x"5f",x"5f",x"00",x"00"),
  1842 => (x"00",x"00",x"00",x"00"),
  1843 => (x"03",x"00",x"03",x"03"),
  1844 => (x"14",x"00",x"00",x"03"),
  1845 => (x"7f",x"14",x"7f",x"7f"),
  1846 => (x"00",x"00",x"14",x"7f"),
  1847 => (x"6b",x"6b",x"2e",x"24"),
  1848 => (x"4c",x"00",x"12",x"3a"),
  1849 => (x"6c",x"18",x"36",x"6a"),
  1850 => (x"30",x"00",x"32",x"56"),
  1851 => (x"77",x"59",x"4f",x"7e"),
  1852 => (x"00",x"40",x"68",x"3a"),
  1853 => (x"03",x"07",x"04",x"00"),
  1854 => (x"00",x"00",x"00",x"00"),
  1855 => (x"63",x"3e",x"1c",x"00"),
  1856 => (x"00",x"00",x"00",x"41"),
  1857 => (x"3e",x"63",x"41",x"00"),
  1858 => (x"08",x"00",x"00",x"1c"),
  1859 => (x"1c",x"1c",x"3e",x"2a"),
  1860 => (x"00",x"08",x"2a",x"3e"),
  1861 => (x"3e",x"3e",x"08",x"08"),
  1862 => (x"00",x"00",x"08",x"08"),
  1863 => (x"60",x"e0",x"80",x"00"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"08",x"08",x"08",x"08"),
  1866 => (x"00",x"00",x"08",x"08"),
  1867 => (x"60",x"60",x"00",x"00"),
  1868 => (x"40",x"00",x"00",x"00"),
  1869 => (x"0c",x"18",x"30",x"60"),
  1870 => (x"00",x"01",x"03",x"06"),
  1871 => (x"4d",x"59",x"7f",x"3e"),
  1872 => (x"00",x"00",x"3e",x"7f"),
  1873 => (x"7f",x"7f",x"06",x"04"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"59",x"71",x"63",x"42"),
  1876 => (x"00",x"00",x"46",x"4f"),
  1877 => (x"49",x"49",x"63",x"22"),
  1878 => (x"18",x"00",x"36",x"7f"),
  1879 => (x"7f",x"13",x"16",x"1c"),
  1880 => (x"00",x"00",x"10",x"7f"),
  1881 => (x"45",x"45",x"67",x"27"),
  1882 => (x"00",x"00",x"39",x"7d"),
  1883 => (x"49",x"4b",x"7e",x"3c"),
  1884 => (x"00",x"00",x"30",x"79"),
  1885 => (x"79",x"71",x"01",x"01"),
  1886 => (x"00",x"00",x"07",x"0f"),
  1887 => (x"49",x"49",x"7f",x"36"),
  1888 => (x"00",x"00",x"36",x"7f"),
  1889 => (x"69",x"49",x"4f",x"06"),
  1890 => (x"00",x"00",x"1e",x"3f"),
  1891 => (x"66",x"66",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"66",x"e6",x"80",x"00"),
  1894 => (x"00",x"00",x"00",x"00"),
  1895 => (x"14",x"14",x"08",x"08"),
  1896 => (x"00",x"00",x"22",x"22"),
  1897 => (x"14",x"14",x"14",x"14"),
  1898 => (x"00",x"00",x"14",x"14"),
  1899 => (x"14",x"14",x"22",x"22"),
  1900 => (x"00",x"00",x"08",x"08"),
  1901 => (x"59",x"51",x"03",x"02"),
  1902 => (x"3e",x"00",x"06",x"0f"),
  1903 => (x"55",x"5d",x"41",x"7f"),
  1904 => (x"00",x"00",x"1e",x"1f"),
  1905 => (x"09",x"09",x"7f",x"7e"),
  1906 => (x"00",x"00",x"7e",x"7f"),
  1907 => (x"49",x"49",x"7f",x"7f"),
  1908 => (x"00",x"00",x"36",x"7f"),
  1909 => (x"41",x"63",x"3e",x"1c"),
  1910 => (x"00",x"00",x"41",x"41"),
  1911 => (x"63",x"41",x"7f",x"7f"),
  1912 => (x"00",x"00",x"1c",x"3e"),
  1913 => (x"49",x"49",x"7f",x"7f"),
  1914 => (x"00",x"00",x"41",x"41"),
  1915 => (x"09",x"09",x"7f",x"7f"),
  1916 => (x"00",x"00",x"01",x"01"),
  1917 => (x"49",x"41",x"7f",x"3e"),
  1918 => (x"00",x"00",x"7a",x"7b"),
  1919 => (x"08",x"08",x"7f",x"7f"),
  1920 => (x"00",x"00",x"7f",x"7f"),
  1921 => (x"7f",x"7f",x"41",x"00"),
  1922 => (x"00",x"00",x"00",x"41"),
  1923 => (x"40",x"40",x"60",x"20"),
  1924 => (x"7f",x"00",x"3f",x"7f"),
  1925 => (x"36",x"1c",x"08",x"7f"),
  1926 => (x"00",x"00",x"41",x"63"),
  1927 => (x"40",x"40",x"7f",x"7f"),
  1928 => (x"7f",x"00",x"40",x"40"),
  1929 => (x"06",x"0c",x"06",x"7f"),
  1930 => (x"7f",x"00",x"7f",x"7f"),
  1931 => (x"18",x"0c",x"06",x"7f"),
  1932 => (x"00",x"00",x"7f",x"7f"),
  1933 => (x"41",x"41",x"7f",x"3e"),
  1934 => (x"00",x"00",x"3e",x"7f"),
  1935 => (x"09",x"09",x"7f",x"7f"),
  1936 => (x"3e",x"00",x"06",x"0f"),
  1937 => (x"7f",x"61",x"41",x"7f"),
  1938 => (x"00",x"00",x"40",x"7e"),
  1939 => (x"19",x"09",x"7f",x"7f"),
  1940 => (x"00",x"00",x"66",x"7f"),
  1941 => (x"59",x"4d",x"6f",x"26"),
  1942 => (x"00",x"00",x"32",x"7b"),
  1943 => (x"7f",x"7f",x"01",x"01"),
  1944 => (x"00",x"00",x"01",x"01"),
  1945 => (x"40",x"40",x"7f",x"3f"),
  1946 => (x"00",x"00",x"3f",x"7f"),
  1947 => (x"70",x"70",x"3f",x"0f"),
  1948 => (x"7f",x"00",x"0f",x"3f"),
  1949 => (x"30",x"18",x"30",x"7f"),
  1950 => (x"41",x"00",x"7f",x"7f"),
  1951 => (x"1c",x"1c",x"36",x"63"),
  1952 => (x"01",x"41",x"63",x"36"),
  1953 => (x"7c",x"7c",x"06",x"03"),
  1954 => (x"61",x"01",x"03",x"06"),
  1955 => (x"47",x"4d",x"59",x"71"),
  1956 => (x"00",x"00",x"41",x"43"),
  1957 => (x"41",x"7f",x"7f",x"00"),
  1958 => (x"01",x"00",x"00",x"41"),
  1959 => (x"18",x"0c",x"06",x"03"),
  1960 => (x"00",x"40",x"60",x"30"),
  1961 => (x"7f",x"41",x"41",x"00"),
  1962 => (x"08",x"00",x"00",x"7f"),
  1963 => (x"06",x"03",x"06",x"0c"),
  1964 => (x"80",x"00",x"08",x"0c"),
  1965 => (x"80",x"80",x"80",x"80"),
  1966 => (x"00",x"00",x"80",x"80"),
  1967 => (x"07",x"03",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"04"),
  1969 => (x"54",x"54",x"74",x"20"),
  1970 => (x"00",x"00",x"78",x"7c"),
  1971 => (x"44",x"44",x"7f",x"7f"),
  1972 => (x"00",x"00",x"38",x"7c"),
  1973 => (x"44",x"44",x"7c",x"38"),
  1974 => (x"00",x"00",x"00",x"44"),
  1975 => (x"44",x"44",x"7c",x"38"),
  1976 => (x"00",x"00",x"7f",x"7f"),
  1977 => (x"54",x"54",x"7c",x"38"),
  1978 => (x"00",x"00",x"18",x"5c"),
  1979 => (x"05",x"7f",x"7e",x"04"),
  1980 => (x"00",x"00",x"00",x"05"),
  1981 => (x"a4",x"a4",x"bc",x"18"),
  1982 => (x"00",x"00",x"7c",x"fc"),
  1983 => (x"04",x"04",x"7f",x"7f"),
  1984 => (x"00",x"00",x"78",x"7c"),
  1985 => (x"7d",x"3d",x"00",x"00"),
  1986 => (x"00",x"00",x"00",x"40"),
  1987 => (x"fd",x"80",x"80",x"80"),
  1988 => (x"00",x"00",x"00",x"7d"),
  1989 => (x"38",x"10",x"7f",x"7f"),
  1990 => (x"00",x"00",x"44",x"6c"),
  1991 => (x"7f",x"3f",x"00",x"00"),
  1992 => (x"7c",x"00",x"00",x"40"),
  1993 => (x"0c",x"18",x"0c",x"7c"),
  1994 => (x"00",x"00",x"78",x"7c"),
  1995 => (x"04",x"04",x"7c",x"7c"),
  1996 => (x"00",x"00",x"78",x"7c"),
  1997 => (x"44",x"44",x"7c",x"38"),
  1998 => (x"00",x"00",x"38",x"7c"),
  1999 => (x"24",x"24",x"fc",x"fc"),
  2000 => (x"00",x"00",x"18",x"3c"),
  2001 => (x"24",x"24",x"3c",x"18"),
  2002 => (x"00",x"00",x"fc",x"fc"),
  2003 => (x"04",x"04",x"7c",x"7c"),
  2004 => (x"00",x"00",x"08",x"0c"),
  2005 => (x"54",x"54",x"5c",x"48"),
  2006 => (x"00",x"00",x"20",x"74"),
  2007 => (x"44",x"7f",x"3f",x"04"),
  2008 => (x"00",x"00",x"00",x"44"),
  2009 => (x"40",x"40",x"7c",x"3c"),
  2010 => (x"00",x"00",x"7c",x"7c"),
  2011 => (x"60",x"60",x"3c",x"1c"),
  2012 => (x"3c",x"00",x"1c",x"3c"),
  2013 => (x"60",x"30",x"60",x"7c"),
  2014 => (x"44",x"00",x"3c",x"7c"),
  2015 => (x"38",x"10",x"38",x"6c"),
  2016 => (x"00",x"00",x"44",x"6c"),
  2017 => (x"60",x"e0",x"bc",x"1c"),
  2018 => (x"00",x"00",x"1c",x"3c"),
  2019 => (x"5c",x"74",x"64",x"44"),
  2020 => (x"00",x"00",x"44",x"4c"),
  2021 => (x"77",x"3e",x"08",x"08"),
  2022 => (x"00",x"00",x"41",x"41"),
  2023 => (x"7f",x"7f",x"00",x"00"),
  2024 => (x"00",x"00",x"00",x"00"),
  2025 => (x"3e",x"77",x"41",x"41"),
  2026 => (x"02",x"00",x"08",x"08"),
  2027 => (x"02",x"03",x"01",x"01"),
  2028 => (x"7f",x"00",x"01",x"02"),
  2029 => (x"7f",x"7f",x"7f",x"7f"),
  2030 => (x"08",x"00",x"7f",x"7f"),
  2031 => (x"3e",x"1c",x"1c",x"08"),
  2032 => (x"7f",x"7f",x"7f",x"3e"),
  2033 => (x"1c",x"3e",x"3e",x"7f"),
  2034 => (x"00",x"08",x"08",x"1c"),
  2035 => (x"7c",x"7c",x"18",x"10"),
  2036 => (x"00",x"00",x"10",x"18"),
  2037 => (x"7c",x"7c",x"30",x"10"),
  2038 => (x"10",x"00",x"10",x"30"),
  2039 => (x"78",x"60",x"60",x"30"),
  2040 => (x"42",x"00",x"06",x"1e"),
  2041 => (x"3c",x"18",x"3c",x"66"),
  2042 => (x"78",x"00",x"42",x"66"),
  2043 => (x"c6",x"c2",x"6a",x"38"),
  2044 => (x"60",x"00",x"38",x"6c"),
  2045 => (x"00",x"60",x"00",x"00"),
  2046 => (x"0e",x"00",x"60",x"00"),
  2047 => (x"5d",x"5c",x"5b",x"5e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

