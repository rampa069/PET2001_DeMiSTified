
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"4c",x"71",x"1e",x"0e"),
     1 => (x"bf",x"d1",x"f4",x"c2"),
     2 => (x"c0",x"4b",x"c0",x"4d"),
     3 => (x"02",x"ab",x"74",x"1e"),
     4 => (x"a6",x"c4",x"87",x"c7"),
     5 => (x"c5",x"78",x"c0",x"48"),
     6 => (x"48",x"a6",x"c4",x"87"),
     7 => (x"66",x"c4",x"78",x"c1"),
     8 => (x"ee",x"49",x"73",x"1e"),
     9 => (x"86",x"c8",x"87",x"df"),
    10 => (x"ef",x"49",x"e0",x"c0"),
    11 => (x"a5",x"c4",x"87",x"ef"),
    12 => (x"f0",x"49",x"6a",x"4a"),
    13 => (x"c6",x"f1",x"87",x"f0"),
    14 => (x"c1",x"85",x"cb",x"87"),
    15 => (x"ab",x"b7",x"c8",x"83"),
    16 => (x"87",x"c7",x"ff",x"04"),
    17 => (x"26",x"4d",x"26",x"26"),
    18 => (x"26",x"4b",x"26",x"4c"),
    19 => (x"4a",x"71",x"1e",x"4f"),
    20 => (x"5a",x"d5",x"f4",x"c2"),
    21 => (x"48",x"d5",x"f4",x"c2"),
    22 => (x"fe",x"49",x"78",x"c7"),
    23 => (x"4f",x"26",x"87",x"dd"),
    24 => (x"71",x"1e",x"73",x"1e"),
    25 => (x"aa",x"b7",x"c0",x"4a"),
    26 => (x"c2",x"87",x"d3",x"03"),
    27 => (x"05",x"bf",x"de",x"cf"),
    28 => (x"4b",x"c1",x"87",x"c4"),
    29 => (x"4b",x"c0",x"87",x"c2"),
    30 => (x"5b",x"e2",x"cf",x"c2"),
    31 => (x"cf",x"c2",x"87",x"c4"),
    32 => (x"cf",x"c2",x"5a",x"e2"),
    33 => (x"c1",x"4a",x"bf",x"de"),
    34 => (x"a2",x"c0",x"c1",x"9a"),
    35 => (x"87",x"e8",x"ec",x"49"),
    36 => (x"cf",x"c2",x"48",x"fc"),
    37 => (x"fe",x"78",x"bf",x"de"),
    38 => (x"71",x"1e",x"87",x"ef"),
    39 => (x"1e",x"66",x"c4",x"4a"),
    40 => (x"f9",x"e9",x"49",x"72"),
    41 => (x"4f",x"26",x"26",x"87"),
    42 => (x"ff",x"4a",x"71",x"1e"),
    43 => (x"ff",x"c3",x"48",x"d4"),
    44 => (x"48",x"d0",x"ff",x"78"),
    45 => (x"ff",x"78",x"e1",x"c0"),
    46 => (x"78",x"c1",x"48",x"d4"),
    47 => (x"31",x"c4",x"49",x"72"),
    48 => (x"d0",x"ff",x"78",x"71"),
    49 => (x"78",x"e0",x"c0",x"48"),
    50 => (x"c2",x"1e",x"4f",x"26"),
    51 => (x"49",x"bf",x"de",x"cf"),
    52 => (x"c2",x"87",x"cc",x"da"),
    53 => (x"e8",x"48",x"c9",x"f4"),
    54 => (x"f4",x"c2",x"78",x"bf"),
    55 => (x"bf",x"ec",x"48",x"c5"),
    56 => (x"c9",x"f4",x"c2",x"78"),
    57 => (x"c3",x"49",x"4a",x"bf"),
    58 => (x"b7",x"c8",x"99",x"ff"),
    59 => (x"71",x"48",x"72",x"2a"),
    60 => (x"d1",x"f4",x"c2",x"b0"),
    61 => (x"0e",x"4f",x"26",x"58"),
    62 => (x"5d",x"5c",x"5b",x"5e"),
    63 => (x"ff",x"4b",x"71",x"0e"),
    64 => (x"f4",x"c2",x"87",x"c8"),
    65 => (x"50",x"c0",x"48",x"c4"),
    66 => (x"ee",x"e5",x"49",x"73"),
    67 => (x"4c",x"49",x"70",x"87"),
    68 => (x"ee",x"cb",x"9c",x"c2"),
    69 => (x"87",x"ce",x"cb",x"49"),
    70 => (x"c2",x"4d",x"49",x"70"),
    71 => (x"bf",x"97",x"c4",x"f4"),
    72 => (x"87",x"e2",x"c1",x"05"),
    73 => (x"c2",x"49",x"66",x"d0"),
    74 => (x"99",x"bf",x"cd",x"f4"),
    75 => (x"d4",x"87",x"d6",x"05"),
    76 => (x"f4",x"c2",x"49",x"66"),
    77 => (x"05",x"99",x"bf",x"c5"),
    78 => (x"49",x"73",x"87",x"cb"),
    79 => (x"70",x"87",x"fc",x"e4"),
    80 => (x"c1",x"c1",x"02",x"98"),
    81 => (x"fe",x"4c",x"c1",x"87"),
    82 => (x"49",x"75",x"87",x"c0"),
    83 => (x"70",x"87",x"e3",x"ca"),
    84 => (x"87",x"c6",x"02",x"98"),
    85 => (x"48",x"c4",x"f4",x"c2"),
    86 => (x"f4",x"c2",x"50",x"c1"),
    87 => (x"05",x"bf",x"97",x"c4"),
    88 => (x"c2",x"87",x"e3",x"c0"),
    89 => (x"49",x"bf",x"cd",x"f4"),
    90 => (x"05",x"99",x"66",x"d0"),
    91 => (x"c2",x"87",x"d6",x"ff"),
    92 => (x"49",x"bf",x"c5",x"f4"),
    93 => (x"05",x"99",x"66",x"d4"),
    94 => (x"73",x"87",x"ca",x"ff"),
    95 => (x"87",x"fb",x"e3",x"49"),
    96 => (x"fe",x"05",x"98",x"70"),
    97 => (x"48",x"74",x"87",x"ff"),
    98 => (x"0e",x"87",x"fa",x"fa"),
    99 => (x"5d",x"5c",x"5b",x"5e"),
   100 => (x"c0",x"86",x"f8",x"0e"),
   101 => (x"bf",x"ec",x"4c",x"4d"),
   102 => (x"48",x"a6",x"c4",x"7e"),
   103 => (x"bf",x"d1",x"f4",x"c2"),
   104 => (x"c0",x"1e",x"c1",x"78"),
   105 => (x"fd",x"49",x"c7",x"1e"),
   106 => (x"86",x"c8",x"87",x"cd"),
   107 => (x"cd",x"02",x"98",x"70"),
   108 => (x"fa",x"49",x"ff",x"87"),
   109 => (x"da",x"c1",x"87",x"ea"),
   110 => (x"87",x"ff",x"e2",x"49"),
   111 => (x"f4",x"c2",x"4d",x"c1"),
   112 => (x"02",x"bf",x"97",x"c4"),
   113 => (x"cf",x"c2",x"87",x"cf"),
   114 => (x"c1",x"49",x"bf",x"d6"),
   115 => (x"da",x"cf",x"c2",x"b9"),
   116 => (x"d3",x"fb",x"71",x"59"),
   117 => (x"c9",x"f4",x"c2",x"87"),
   118 => (x"cf",x"c2",x"4b",x"bf"),
   119 => (x"c0",x"05",x"bf",x"de"),
   120 => (x"fd",x"c3",x"87",x"e9"),
   121 => (x"87",x"d3",x"e2",x"49"),
   122 => (x"e2",x"49",x"fa",x"c3"),
   123 => (x"49",x"73",x"87",x"cd"),
   124 => (x"71",x"99",x"ff",x"c3"),
   125 => (x"fa",x"49",x"c0",x"1e"),
   126 => (x"49",x"73",x"87",x"e0"),
   127 => (x"71",x"29",x"b7",x"c8"),
   128 => (x"fa",x"49",x"c1",x"1e"),
   129 => (x"86",x"c8",x"87",x"d4"),
   130 => (x"c2",x"87",x"f5",x"c5"),
   131 => (x"4b",x"bf",x"cd",x"f4"),
   132 => (x"87",x"dd",x"02",x"9b"),
   133 => (x"bf",x"da",x"cf",x"c2"),
   134 => (x"87",x"d6",x"c7",x"49"),
   135 => (x"c4",x"05",x"98",x"70"),
   136 => (x"d2",x"4b",x"c0",x"87"),
   137 => (x"49",x"e0",x"c2",x"87"),
   138 => (x"c2",x"87",x"fb",x"c6"),
   139 => (x"c6",x"58",x"de",x"cf"),
   140 => (x"da",x"cf",x"c2",x"87"),
   141 => (x"73",x"78",x"c0",x"48"),
   142 => (x"05",x"99",x"c2",x"49"),
   143 => (x"eb",x"c3",x"87",x"cd"),
   144 => (x"87",x"f7",x"e0",x"49"),
   145 => (x"99",x"c2",x"49",x"70"),
   146 => (x"fb",x"87",x"c2",x"02"),
   147 => (x"c1",x"49",x"73",x"4c"),
   148 => (x"87",x"cd",x"05",x"99"),
   149 => (x"e0",x"49",x"f4",x"c3"),
   150 => (x"49",x"70",x"87",x"e1"),
   151 => (x"c2",x"02",x"99",x"c2"),
   152 => (x"73",x"4c",x"fa",x"87"),
   153 => (x"05",x"99",x"c8",x"49"),
   154 => (x"f5",x"c3",x"87",x"cd"),
   155 => (x"87",x"cb",x"e0",x"49"),
   156 => (x"99",x"c2",x"49",x"70"),
   157 => (x"c2",x"87",x"d5",x"02"),
   158 => (x"02",x"bf",x"d5",x"f4"),
   159 => (x"c1",x"48",x"87",x"ca"),
   160 => (x"d9",x"f4",x"c2",x"88"),
   161 => (x"87",x"c2",x"c0",x"58"),
   162 => (x"4d",x"c1",x"4c",x"ff"),
   163 => (x"99",x"c4",x"49",x"73"),
   164 => (x"c3",x"87",x"ce",x"05"),
   165 => (x"df",x"ff",x"49",x"f2"),
   166 => (x"49",x"70",x"87",x"e1"),
   167 => (x"dc",x"02",x"99",x"c2"),
   168 => (x"d5",x"f4",x"c2",x"87"),
   169 => (x"c7",x"48",x"7e",x"bf"),
   170 => (x"c0",x"03",x"a8",x"b7"),
   171 => (x"48",x"6e",x"87",x"cb"),
   172 => (x"f4",x"c2",x"80",x"c1"),
   173 => (x"c2",x"c0",x"58",x"d9"),
   174 => (x"c1",x"4c",x"fe",x"87"),
   175 => (x"49",x"fd",x"c3",x"4d"),
   176 => (x"87",x"f7",x"de",x"ff"),
   177 => (x"99",x"c2",x"49",x"70"),
   178 => (x"c2",x"87",x"d5",x"02"),
   179 => (x"02",x"bf",x"d5",x"f4"),
   180 => (x"c2",x"87",x"c9",x"c0"),
   181 => (x"c0",x"48",x"d5",x"f4"),
   182 => (x"87",x"c2",x"c0",x"78"),
   183 => (x"4d",x"c1",x"4c",x"fd"),
   184 => (x"ff",x"49",x"fa",x"c3"),
   185 => (x"70",x"87",x"d4",x"de"),
   186 => (x"02",x"99",x"c2",x"49"),
   187 => (x"c2",x"87",x"d9",x"c0"),
   188 => (x"48",x"bf",x"d5",x"f4"),
   189 => (x"03",x"a8",x"b7",x"c7"),
   190 => (x"c2",x"87",x"c9",x"c0"),
   191 => (x"c7",x"48",x"d5",x"f4"),
   192 => (x"87",x"c2",x"c0",x"78"),
   193 => (x"4d",x"c1",x"4c",x"fc"),
   194 => (x"03",x"ac",x"b7",x"c0"),
   195 => (x"c4",x"87",x"d3",x"c0"),
   196 => (x"d8",x"c1",x"48",x"66"),
   197 => (x"6e",x"7e",x"70",x"80"),
   198 => (x"c5",x"c0",x"02",x"bf"),
   199 => (x"49",x"74",x"4b",x"87"),
   200 => (x"1e",x"c0",x"0f",x"73"),
   201 => (x"c1",x"1e",x"f0",x"c3"),
   202 => (x"ca",x"f7",x"49",x"da"),
   203 => (x"70",x"86",x"c8",x"87"),
   204 => (x"d8",x"c0",x"02",x"98"),
   205 => (x"d5",x"f4",x"c2",x"87"),
   206 => (x"49",x"6e",x"7e",x"bf"),
   207 => (x"66",x"c4",x"91",x"cb"),
   208 => (x"6a",x"82",x"71",x"4a"),
   209 => (x"87",x"c5",x"c0",x"02"),
   210 => (x"73",x"49",x"6e",x"4b"),
   211 => (x"02",x"9d",x"75",x"0f"),
   212 => (x"c2",x"87",x"c8",x"c0"),
   213 => (x"49",x"bf",x"d5",x"f4"),
   214 => (x"c2",x"87",x"e0",x"f2"),
   215 => (x"02",x"bf",x"e2",x"cf"),
   216 => (x"49",x"87",x"dd",x"c0"),
   217 => (x"70",x"87",x"cb",x"c2"),
   218 => (x"d3",x"c0",x"02",x"98"),
   219 => (x"d5",x"f4",x"c2",x"87"),
   220 => (x"c6",x"f2",x"49",x"bf"),
   221 => (x"f3",x"49",x"c0",x"87"),
   222 => (x"cf",x"c2",x"87",x"e6"),
   223 => (x"78",x"c0",x"48",x"e2"),
   224 => (x"c0",x"f3",x"8e",x"f8"),
   225 => (x"5b",x"5e",x"0e",x"87"),
   226 => (x"1e",x"0e",x"5d",x"5c"),
   227 => (x"f4",x"c2",x"4c",x"71"),
   228 => (x"c1",x"49",x"bf",x"d1"),
   229 => (x"c1",x"4d",x"a1",x"cd"),
   230 => (x"7e",x"69",x"81",x"d1"),
   231 => (x"cf",x"02",x"9c",x"74"),
   232 => (x"4b",x"a5",x"c4",x"87"),
   233 => (x"f4",x"c2",x"7b",x"74"),
   234 => (x"f2",x"49",x"bf",x"d1"),
   235 => (x"7b",x"6e",x"87",x"df"),
   236 => (x"c4",x"05",x"9c",x"74"),
   237 => (x"c2",x"4b",x"c0",x"87"),
   238 => (x"73",x"4b",x"c1",x"87"),
   239 => (x"87",x"e0",x"f2",x"49"),
   240 => (x"c7",x"02",x"66",x"d4"),
   241 => (x"87",x"de",x"49",x"87"),
   242 => (x"87",x"c2",x"4a",x"70"),
   243 => (x"cf",x"c2",x"4a",x"c0"),
   244 => (x"f1",x"26",x"5a",x"e6"),
   245 => (x"00",x"00",x"87",x"ef"),
   246 => (x"00",x"00",x"00",x"00"),
   247 => (x"00",x"00",x"00",x"00"),
   248 => (x"00",x"00",x"00",x"00"),
   249 => (x"71",x"1e",x"00",x"00"),
   250 => (x"bf",x"c8",x"ff",x"4a"),
   251 => (x"48",x"a1",x"72",x"49"),
   252 => (x"ff",x"1e",x"4f",x"26"),
   253 => (x"fe",x"89",x"bf",x"c8"),
   254 => (x"c0",x"c0",x"c0",x"c0"),
   255 => (x"c4",x"01",x"a9",x"c0"),
   256 => (x"c2",x"4a",x"c0",x"87"),
   257 => (x"72",x"4a",x"c1",x"87"),
   258 => (x"1e",x"4f",x"26",x"48"),
   259 => (x"87",x"db",x"d2",x"ff"),
   260 => (x"c2",x"49",x"66",x"c4"),
   261 => (x"cd",x"02",x"99",x"c0"),
   262 => (x"1e",x"e0",x"c3",x"87"),
   263 => (x"49",x"e6",x"f3",x"c2"),
   264 => (x"87",x"ea",x"d3",x"ff"),
   265 => (x"66",x"c4",x"86",x"c4"),
   266 => (x"99",x"c0",x"c4",x"49"),
   267 => (x"c3",x"87",x"cd",x"02"),
   268 => (x"f3",x"c2",x"1e",x"f0"),
   269 => (x"d3",x"ff",x"49",x"e6"),
   270 => (x"86",x"c4",x"87",x"d4"),
   271 => (x"c1",x"49",x"66",x"c4"),
   272 => (x"1e",x"71",x"99",x"ff"),
   273 => (x"49",x"e6",x"f3",x"c2"),
   274 => (x"87",x"c2",x"d3",x"ff"),
   275 => (x"87",x"d3",x"d1",x"ff"),
   276 => (x"0e",x"4f",x"26",x"26"),
   277 => (x"5d",x"5c",x"5b",x"5e"),
   278 => (x"86",x"dc",x"ff",x"0e"),
   279 => (x"f4",x"c2",x"7e",x"c0"),
   280 => (x"c2",x"49",x"bf",x"dd"),
   281 => (x"72",x"1e",x"71",x"81"),
   282 => (x"fd",x"4a",x"c6",x"1e"),
   283 => (x"71",x"87",x"fc",x"f1"),
   284 => (x"26",x"4a",x"26",x"48"),
   285 => (x"58",x"a6",x"c8",x"49"),
   286 => (x"bf",x"dd",x"f4",x"c2"),
   287 => (x"71",x"81",x"c4",x"49"),
   288 => (x"c6",x"1e",x"72",x"1e"),
   289 => (x"e2",x"f1",x"fd",x"4a"),
   290 => (x"26",x"48",x"71",x"87"),
   291 => (x"cc",x"49",x"26",x"4a"),
   292 => (x"dc",x"c2",x"58",x"a6"),
   293 => (x"fd",x"49",x"bf",x"f9"),
   294 => (x"98",x"70",x"87",x"d8"),
   295 => (x"87",x"ce",x"ca",x"02"),
   296 => (x"fd",x"49",x"e0",x"c0"),
   297 => (x"49",x"70",x"87",x"c0"),
   298 => (x"59",x"fd",x"dc",x"c2"),
   299 => (x"49",x"74",x"4c",x"c0"),
   300 => (x"d0",x"fe",x"91",x"c4"),
   301 => (x"74",x"4a",x"69",x"81"),
   302 => (x"dd",x"f4",x"c2",x"49"),
   303 => (x"91",x"c4",x"81",x"bf"),
   304 => (x"81",x"ed",x"f4",x"c2"),
   305 => (x"02",x"9a",x"79",x"72"),
   306 => (x"49",x"72",x"87",x"d2"),
   307 => (x"9a",x"71",x"89",x"c1"),
   308 => (x"80",x"c1",x"48",x"6e"),
   309 => (x"9a",x"72",x"7e",x"70"),
   310 => (x"87",x"ee",x"ff",x"05"),
   311 => (x"b7",x"c2",x"84",x"c1"),
   312 => (x"c9",x"ff",x"04",x"ac"),
   313 => (x"c0",x"48",x"6e",x"87"),
   314 => (x"04",x"a8",x"b7",x"fc"),
   315 => (x"c0",x"87",x"ff",x"c8"),
   316 => (x"c4",x"4a",x"74",x"4c"),
   317 => (x"92",x"c4",x"82",x"66"),
   318 => (x"82",x"ed",x"f4",x"c2"),
   319 => (x"66",x"c8",x"49",x"74"),
   320 => (x"c2",x"91",x"c4",x"81"),
   321 => (x"6a",x"81",x"ed",x"f4"),
   322 => (x"72",x"49",x"69",x"4a"),
   323 => (x"c2",x"4b",x"74",x"b9"),
   324 => (x"83",x"bf",x"dd",x"f4"),
   325 => (x"f4",x"c2",x"93",x"c4"),
   326 => (x"ba",x"6b",x"83",x"ed"),
   327 => (x"98",x"71",x"48",x"72"),
   328 => (x"74",x"58",x"a6",x"d0"),
   329 => (x"dd",x"f4",x"c2",x"49"),
   330 => (x"91",x"c4",x"81",x"bf"),
   331 => (x"81",x"ed",x"f4",x"c2"),
   332 => (x"a6",x"d0",x"7e",x"69"),
   333 => (x"cc",x"78",x"c0",x"48"),
   334 => (x"29",x"df",x"49",x"66"),
   335 => (x"87",x"c0",x"c7",x"02"),
   336 => (x"e0",x"c0",x"4a",x"74"),
   337 => (x"82",x"66",x"d0",x"92"),
   338 => (x"72",x"48",x"ff",x"c0"),
   339 => (x"d4",x"4a",x"70",x"88"),
   340 => (x"78",x"c0",x"48",x"a6"),
   341 => (x"78",x"c0",x"80",x"c4"),
   342 => (x"29",x"df",x"49",x"6e"),
   343 => (x"59",x"a6",x"e0",x"c0"),
   344 => (x"48",x"d9",x"f4",x"c2"),
   345 => (x"49",x"72",x"78",x"c1"),
   346 => (x"2a",x"b7",x"31",x"c3"),
   347 => (x"ff",x"c0",x"b1",x"72"),
   348 => (x"c2",x"91",x"c4",x"99"),
   349 => (x"71",x"4d",x"d0",x"de"),
   350 => (x"49",x"4b",x"6d",x"85"),
   351 => (x"99",x"c0",x"c0",x"c4"),
   352 => (x"87",x"f3",x"c0",x"02"),
   353 => (x"c8",x"02",x"66",x"dc"),
   354 => (x"c0",x"80",x"c8",x"87"),
   355 => (x"ef",x"c5",x"78",x"40"),
   356 => (x"e1",x"f4",x"c2",x"87"),
   357 => (x"c2",x"78",x"c1",x"48"),
   358 => (x"05",x"bf",x"e5",x"f4"),
   359 => (x"c1",x"87",x"e1",x"c5"),
   360 => (x"a0",x"f8",x"1e",x"d8"),
   361 => (x"87",x"e3",x"f9",x"49"),
   362 => (x"c2",x"1e",x"d8",x"c5"),
   363 => (x"f9",x"49",x"d9",x"f4"),
   364 => (x"86",x"c8",x"87",x"d9"),
   365 => (x"dc",x"87",x"c9",x"c5"),
   366 => (x"87",x"d8",x"02",x"66"),
   367 => (x"c0",x"c2",x"49",x"73"),
   368 => (x"c0",x"02",x"99",x"c0"),
   369 => (x"b7",x"d0",x"87",x"c3"),
   370 => (x"fd",x"48",x"6d",x"2b"),
   371 => (x"70",x"98",x"ff",x"ff"),
   372 => (x"87",x"fa",x"c0",x"7d"),
   373 => (x"bf",x"e1",x"f4",x"c2"),
   374 => (x"87",x"f2",x"c0",x"02"),
   375 => (x"b7",x"d0",x"48",x"73"),
   376 => (x"a6",x"e4",x"c0",x"28"),
   377 => (x"02",x"98",x"70",x"58"),
   378 => (x"c2",x"87",x"e3",x"c0"),
   379 => (x"49",x"bf",x"e9",x"f4"),
   380 => (x"99",x"c0",x"e0",x"c0"),
   381 => (x"87",x"ca",x"c0",x"02"),
   382 => (x"e0",x"c0",x"49",x"70"),
   383 => (x"c0",x"02",x"99",x"c0"),
   384 => (x"48",x"6d",x"87",x"cc"),
   385 => (x"b0",x"c0",x"c0",x"c2"),
   386 => (x"e0",x"c0",x"7d",x"70"),
   387 => (x"49",x"73",x"4b",x"66"),
   388 => (x"99",x"c0",x"c0",x"c8"),
   389 => (x"87",x"c7",x"c2",x"02"),
   390 => (x"bf",x"e9",x"f4",x"c2"),
   391 => (x"9a",x"c0",x"cc",x"4a"),
   392 => (x"87",x"cf",x"c0",x"02"),
   393 => (x"02",x"8a",x"c0",x"c4"),
   394 => (x"8a",x"87",x"d8",x"c0"),
   395 => (x"87",x"f9",x"c0",x"02"),
   396 => (x"73",x"87",x"dd",x"c1"),
   397 => (x"99",x"ff",x"c3",x"49"),
   398 => (x"de",x"c2",x"91",x"c2"),
   399 => (x"4b",x"11",x"81",x"c4"),
   400 => (x"73",x"87",x"dc",x"c1"),
   401 => (x"99",x"ff",x"c3",x"49"),
   402 => (x"de",x"c2",x"91",x"c2"),
   403 => (x"81",x"c1",x"81",x"c4"),
   404 => (x"66",x"dc",x"4b",x"11"),
   405 => (x"87",x"c8",x"c0",x"02"),
   406 => (x"d2",x"48",x"a6",x"d8"),
   407 => (x"87",x"ff",x"c0",x"78"),
   408 => (x"c4",x"48",x"a6",x"d4"),
   409 => (x"f6",x"c0",x"78",x"d2"),
   410 => (x"c3",x"49",x"73",x"87"),
   411 => (x"91",x"c2",x"99",x"ff"),
   412 => (x"81",x"c4",x"de",x"c2"),
   413 => (x"4b",x"11",x"81",x"c1"),
   414 => (x"c0",x"02",x"66",x"dc"),
   415 => (x"a6",x"d8",x"87",x"c9"),
   416 => (x"78",x"d9",x"c1",x"48"),
   417 => (x"d4",x"87",x"d8",x"c0"),
   418 => (x"d9",x"c5",x"48",x"a6"),
   419 => (x"87",x"cf",x"c0",x"78"),
   420 => (x"ff",x"c3",x"49",x"73"),
   421 => (x"c2",x"91",x"c2",x"99"),
   422 => (x"c1",x"81",x"c4",x"de"),
   423 => (x"dc",x"4b",x"11",x"81"),
   424 => (x"dc",x"c0",x"02",x"66"),
   425 => (x"ff",x"49",x"73",x"87"),
   426 => (x"c0",x"fc",x"c7",x"b9"),
   427 => (x"c2",x"48",x"71",x"99"),
   428 => (x"98",x"bf",x"e9",x"f4"),
   429 => (x"58",x"ed",x"f4",x"c2"),
   430 => (x"c4",x"9b",x"ff",x"c3"),
   431 => (x"d4",x"c0",x"b3",x"c0"),
   432 => (x"c7",x"49",x"73",x"87"),
   433 => (x"71",x"99",x"c0",x"fc"),
   434 => (x"e9",x"f4",x"c2",x"48"),
   435 => (x"f4",x"c2",x"b0",x"bf"),
   436 => (x"ff",x"c3",x"58",x"ed"),
   437 => (x"02",x"66",x"d4",x"9b"),
   438 => (x"1e",x"87",x"ca",x"c0"),
   439 => (x"49",x"d9",x"f4",x"c2"),
   440 => (x"c4",x"87",x"e8",x"f4"),
   441 => (x"c2",x"1e",x"73",x"86"),
   442 => (x"f4",x"49",x"d9",x"f4"),
   443 => (x"86",x"c4",x"87",x"dd"),
   444 => (x"c0",x"02",x"66",x"d8"),
   445 => (x"c2",x"1e",x"87",x"ca"),
   446 => (x"f4",x"49",x"d9",x"f4"),
   447 => (x"86",x"c4",x"87",x"cd"),
   448 => (x"c1",x"48",x"66",x"cc"),
   449 => (x"58",x"a6",x"d0",x"30"),
   450 => (x"30",x"c1",x"48",x"6e"),
   451 => (x"66",x"d0",x"7e",x"70"),
   452 => (x"d4",x"80",x"c1",x"48"),
   453 => (x"e0",x"c0",x"58",x"a6"),
   454 => (x"f8",x"04",x"a8",x"b7"),
   455 => (x"84",x"c1",x"87",x"d9"),
   456 => (x"04",x"ac",x"b7",x"c2"),
   457 => (x"c2",x"87",x"ca",x"f7"),
   458 => (x"c4",x"48",x"dd",x"f4"),
   459 => (x"dc",x"ff",x"78",x"66"),
   460 => (x"26",x"4d",x"26",x"8e"),
   461 => (x"26",x"4b",x"26",x"4c"),
   462 => (x"00",x"00",x"00",x"4f"),
   463 => (x"4a",x"c0",x"1e",x"00"),
   464 => (x"91",x"c4",x"49",x"72"),
   465 => (x"81",x"ed",x"f4",x"c2"),
   466 => (x"82",x"c1",x"79",x"ff"),
   467 => (x"04",x"aa",x"b7",x"c6"),
   468 => (x"f4",x"c2",x"87",x"ee"),
   469 => (x"40",x"c0",x"48",x"dd"),
   470 => (x"c0",x"80",x"c8",x"78"),
   471 => (x"1e",x"4f",x"26",x"78"),
   472 => (x"4b",x"71",x"1e",x"73"),
   473 => (x"bf",x"c0",x"de",x"c2"),
   474 => (x"c2",x"87",x"c9",x"05"),
   475 => (x"c1",x"48",x"c0",x"de"),
   476 => (x"87",x"c9",x"ff",x"78"),
   477 => (x"73",x"87",x"dc",x"f3"),
   478 => (x"fb",x"c7",x"ff",x"49"),
   479 => (x"87",x"f5",x"fe",x"87"),
   480 => (x"00",x"00",x"00",x"00"),
   481 => (x"f5",x"f2",x"eb",x"f4"),
   482 => (x"0c",x"04",x"06",x"05"),
   483 => (x"0a",x"83",x"0b",x"03"),
   484 => (x"00",x"fc",x"00",x"66"),
   485 => (x"00",x"da",x"00",x"5a"),
   486 => (x"08",x"94",x"80",x"00"),
   487 => (x"00",x"78",x"80",x"05"),
   488 => (x"00",x"01",x"80",x"02"),
   489 => (x"00",x"09",x"80",x"03"),
   490 => (x"00",x"00",x"80",x"04"),
   491 => (x"08",x"91",x"80",x"01"),
   492 => (x"00",x"04",x"00",x"26"),
   493 => (x"00",x"00",x"00",x"1d"),
   494 => (x"00",x"00",x"00",x"1c"),
   495 => (x"00",x"0c",x"00",x"25"),
   496 => (x"00",x"00",x"00",x"1a"),
   497 => (x"00",x"00",x"00",x"1b"),
   498 => (x"00",x"00",x"00",x"24"),
   499 => (x"00",x"00",x"01",x"12"),
   500 => (x"00",x"03",x"00",x"2e"),
   501 => (x"00",x"00",x"00",x"2d"),
   502 => (x"00",x"00",x"00",x"23"),
   503 => (x"00",x"0b",x"00",x"36"),
   504 => (x"00",x"00",x"00",x"21"),
   505 => (x"00",x"00",x"00",x"2b"),
   506 => (x"00",x"00",x"00",x"2c"),
   507 => (x"00",x"00",x"00",x"22"),
   508 => (x"00",x"6c",x"00",x"3d"),
   509 => (x"00",x"00",x"00",x"35"),
   510 => (x"00",x"00",x"00",x"34"),
   511 => (x"00",x"75",x"00",x"3e"),
   512 => (x"00",x"00",x"00",x"32"),
   513 => (x"00",x"00",x"00",x"33"),
   514 => (x"00",x"6b",x"00",x"3c"),
   515 => (x"00",x"00",x"00",x"2a"),
   516 => (x"00",x"01",x"00",x"46"),
   517 => (x"00",x"73",x"00",x"43"),
   518 => (x"00",x"69",x"00",x"3b"),
   519 => (x"00",x"09",x"00",x"45"),
   520 => (x"00",x"70",x"00",x"3a"),
   521 => (x"00",x"72",x"00",x"42"),
   522 => (x"00",x"74",x"00",x"44"),
   523 => (x"00",x"00",x"00",x"31"),
   524 => (x"00",x"00",x"00",x"55"),
   525 => (x"00",x"7c",x"00",x"4d"),
   526 => (x"00",x"7a",x"00",x"4b"),
   527 => (x"00",x"00",x"00",x"7b"),
   528 => (x"00",x"71",x"00",x"49"),
   529 => (x"00",x"84",x"00",x"4c"),
   530 => (x"00",x"77",x"00",x"54"),
   531 => (x"00",x"00",x"00",x"41"),
   532 => (x"00",x"00",x"00",x"61"),
   533 => (x"00",x"7c",x"00",x"5b"),
   534 => (x"00",x"00",x"00",x"52"),
   535 => (x"00",x"00",x"00",x"f1"),
   536 => (x"00",x"00",x"02",x"59"),
   537 => (x"00",x"5d",x"00",x"0e"),
   538 => (x"00",x"00",x"00",x"5d"),
   539 => (x"00",x"79",x"00",x"4a"),
   540 => (x"00",x"05",x"00",x"16"),
   541 => (x"00",x"07",x"00",x"76"),
   542 => (x"00",x"0d",x"00",x"0d"),
   543 => (x"00",x"06",x"00",x"1e"),
   544 => (x"00",x"00",x"00",x"29"),
   545 => (x"00",x"00",x"04",x"14"),
   546 => (x"00",x"00",x"00",x"15"),
   547 => (x"00",x"00",x"40",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

