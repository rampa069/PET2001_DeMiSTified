
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"74",x"1e",x"c0",x"4b"),
     1 => (x"87",x"c7",x"02",x"ab"),
     2 => (x"c0",x"48",x"a6",x"c4"),
     3 => (x"c4",x"87",x"c5",x"78"),
     4 => (x"78",x"c1",x"48",x"a6"),
     5 => (x"73",x"1e",x"66",x"c4"),
     6 => (x"87",x"df",x"ee",x"49"),
     7 => (x"e0",x"c0",x"86",x"c8"),
     8 => (x"87",x"ef",x"ef",x"49"),
     9 => (x"6a",x"4a",x"a5",x"c4"),
    10 => (x"87",x"f0",x"f0",x"49"),
    11 => (x"cb",x"87",x"c6",x"f1"),
    12 => (x"c8",x"83",x"c1",x"85"),
    13 => (x"ff",x"04",x"ab",x"b7"),
    14 => (x"26",x"26",x"87",x"c7"),
    15 => (x"26",x"4c",x"26",x"4d"),
    16 => (x"1e",x"4f",x"26",x"4b"),
    17 => (x"f4",x"c2",x"4a",x"71"),
    18 => (x"f4",x"c2",x"5a",x"cd"),
    19 => (x"78",x"c7",x"48",x"cd"),
    20 => (x"87",x"dd",x"fe",x"49"),
    21 => (x"73",x"1e",x"4f",x"26"),
    22 => (x"c0",x"4a",x"71",x"1e"),
    23 => (x"d3",x"03",x"aa",x"b7"),
    24 => (x"d3",x"cf",x"c2",x"87"),
    25 => (x"87",x"c4",x"05",x"bf"),
    26 => (x"87",x"c2",x"4b",x"c1"),
    27 => (x"cf",x"c2",x"4b",x"c0"),
    28 => (x"87",x"c4",x"5b",x"d7"),
    29 => (x"5a",x"d7",x"cf",x"c2"),
    30 => (x"bf",x"d3",x"cf",x"c2"),
    31 => (x"c1",x"9a",x"c1",x"4a"),
    32 => (x"ec",x"49",x"a2",x"c0"),
    33 => (x"48",x"fc",x"87",x"e8"),
    34 => (x"bf",x"d3",x"cf",x"c2"),
    35 => (x"87",x"ef",x"fe",x"78"),
    36 => (x"c4",x"4a",x"71",x"1e"),
    37 => (x"49",x"72",x"1e",x"66"),
    38 => (x"26",x"87",x"f9",x"ea"),
    39 => (x"71",x"1e",x"4f",x"26"),
    40 => (x"48",x"d4",x"ff",x"4a"),
    41 => (x"ff",x"78",x"ff",x"c3"),
    42 => (x"e1",x"c0",x"48",x"d0"),
    43 => (x"48",x"d4",x"ff",x"78"),
    44 => (x"49",x"72",x"78",x"c1"),
    45 => (x"78",x"71",x"31",x"c4"),
    46 => (x"c0",x"48",x"d0",x"ff"),
    47 => (x"4f",x"26",x"78",x"e0"),
    48 => (x"d3",x"cf",x"c2",x"1e"),
    49 => (x"cb",x"da",x"49",x"bf"),
    50 => (x"c1",x"f4",x"c2",x"87"),
    51 => (x"78",x"bf",x"e8",x"48"),
    52 => (x"48",x"fd",x"f3",x"c2"),
    53 => (x"c2",x"78",x"bf",x"ec"),
    54 => (x"4a",x"bf",x"c1",x"f4"),
    55 => (x"99",x"ff",x"c3",x"49"),
    56 => (x"72",x"2a",x"b7",x"c8"),
    57 => (x"c2",x"b0",x"71",x"48"),
    58 => (x"26",x"58",x"c9",x"f4"),
    59 => (x"5b",x"5e",x"0e",x"4f"),
    60 => (x"71",x"0e",x"5d",x"5c"),
    61 => (x"87",x"c8",x"ff",x"4b"),
    62 => (x"48",x"fc",x"f3",x"c2"),
    63 => (x"49",x"73",x"50",x"c0"),
    64 => (x"70",x"87",x"ee",x"e6"),
    65 => (x"9c",x"c2",x"4c",x"49"),
    66 => (x"cb",x"49",x"ee",x"cb"),
    67 => (x"49",x"70",x"87",x"cd"),
    68 => (x"fc",x"f3",x"c2",x"4d"),
    69 => (x"c1",x"05",x"bf",x"97"),
    70 => (x"66",x"d0",x"87",x"e2"),
    71 => (x"c5",x"f4",x"c2",x"49"),
    72 => (x"d6",x"05",x"99",x"bf"),
    73 => (x"49",x"66",x"d4",x"87"),
    74 => (x"bf",x"fd",x"f3",x"c2"),
    75 => (x"87",x"cb",x"05",x"99"),
    76 => (x"fc",x"e5",x"49",x"73"),
    77 => (x"02",x"98",x"70",x"87"),
    78 => (x"c1",x"87",x"c1",x"c1"),
    79 => (x"87",x"c0",x"fe",x"4c"),
    80 => (x"e2",x"ca",x"49",x"75"),
    81 => (x"02",x"98",x"70",x"87"),
    82 => (x"f3",x"c2",x"87",x"c6"),
    83 => (x"50",x"c1",x"48",x"fc"),
    84 => (x"97",x"fc",x"f3",x"c2"),
    85 => (x"e3",x"c0",x"05",x"bf"),
    86 => (x"c5",x"f4",x"c2",x"87"),
    87 => (x"66",x"d0",x"49",x"bf"),
    88 => (x"d6",x"ff",x"05",x"99"),
    89 => (x"fd",x"f3",x"c2",x"87"),
    90 => (x"66",x"d4",x"49",x"bf"),
    91 => (x"ca",x"ff",x"05",x"99"),
    92 => (x"e4",x"49",x"73",x"87"),
    93 => (x"98",x"70",x"87",x"fb"),
    94 => (x"87",x"ff",x"fe",x"05"),
    95 => (x"fa",x"fa",x"48",x"74"),
    96 => (x"5b",x"5e",x"0e",x"87"),
    97 => (x"f8",x"0e",x"5d",x"5c"),
    98 => (x"4c",x"4d",x"c0",x"86"),
    99 => (x"c4",x"7e",x"bf",x"ec"),
   100 => (x"f4",x"c2",x"48",x"a6"),
   101 => (x"c1",x"78",x"bf",x"c9"),
   102 => (x"c7",x"1e",x"c0",x"1e"),
   103 => (x"87",x"cd",x"fd",x"49"),
   104 => (x"98",x"70",x"86",x"c8"),
   105 => (x"ff",x"87",x"cd",x"02"),
   106 => (x"87",x"ea",x"fa",x"49"),
   107 => (x"e3",x"49",x"da",x"c1"),
   108 => (x"4d",x"c1",x"87",x"ff"),
   109 => (x"97",x"fc",x"f3",x"c2"),
   110 => (x"87",x"cf",x"02",x"bf"),
   111 => (x"bf",x"cb",x"cf",x"c2"),
   112 => (x"c2",x"b9",x"c1",x"49"),
   113 => (x"71",x"59",x"cf",x"cf"),
   114 => (x"c2",x"87",x"d3",x"fb"),
   115 => (x"4b",x"bf",x"c1",x"f4"),
   116 => (x"bf",x"d3",x"cf",x"c2"),
   117 => (x"87",x"e9",x"c0",x"05"),
   118 => (x"e3",x"49",x"fd",x"c3"),
   119 => (x"fa",x"c3",x"87",x"d3"),
   120 => (x"87",x"cd",x"e3",x"49"),
   121 => (x"ff",x"c3",x"49",x"73"),
   122 => (x"c0",x"1e",x"71",x"99"),
   123 => (x"87",x"e0",x"fa",x"49"),
   124 => (x"b7",x"c8",x"49",x"73"),
   125 => (x"c1",x"1e",x"71",x"29"),
   126 => (x"87",x"d4",x"fa",x"49"),
   127 => (x"f4",x"c5",x"86",x"c8"),
   128 => (x"c5",x"f4",x"c2",x"87"),
   129 => (x"02",x"9b",x"4b",x"bf"),
   130 => (x"cf",x"c2",x"87",x"dd"),
   131 => (x"c7",x"49",x"bf",x"cf"),
   132 => (x"98",x"70",x"87",x"d5"),
   133 => (x"c0",x"87",x"c4",x"05"),
   134 => (x"c2",x"87",x"d2",x"4b"),
   135 => (x"fa",x"c6",x"49",x"e0"),
   136 => (x"d3",x"cf",x"c2",x"87"),
   137 => (x"c2",x"87",x"c6",x"58"),
   138 => (x"c0",x"48",x"cf",x"cf"),
   139 => (x"c2",x"49",x"73",x"78"),
   140 => (x"87",x"cd",x"05",x"99"),
   141 => (x"e1",x"49",x"eb",x"c3"),
   142 => (x"49",x"70",x"87",x"f7"),
   143 => (x"c2",x"02",x"99",x"c2"),
   144 => (x"73",x"4c",x"fb",x"87"),
   145 => (x"05",x"99",x"c1",x"49"),
   146 => (x"f4",x"c3",x"87",x"cd"),
   147 => (x"87",x"e1",x"e1",x"49"),
   148 => (x"99",x"c2",x"49",x"70"),
   149 => (x"fa",x"87",x"c2",x"02"),
   150 => (x"c8",x"49",x"73",x"4c"),
   151 => (x"87",x"cd",x"05",x"99"),
   152 => (x"e1",x"49",x"f5",x"c3"),
   153 => (x"49",x"70",x"87",x"cb"),
   154 => (x"d5",x"02",x"99",x"c2"),
   155 => (x"cd",x"f4",x"c2",x"87"),
   156 => (x"87",x"ca",x"02",x"bf"),
   157 => (x"c2",x"88",x"c1",x"48"),
   158 => (x"c0",x"58",x"d1",x"f4"),
   159 => (x"4c",x"ff",x"87",x"c2"),
   160 => (x"49",x"73",x"4d",x"c1"),
   161 => (x"cd",x"05",x"99",x"c4"),
   162 => (x"49",x"f2",x"c3",x"87"),
   163 => (x"70",x"87",x"e2",x"e0"),
   164 => (x"02",x"99",x"c2",x"49"),
   165 => (x"f4",x"c2",x"87",x"dc"),
   166 => (x"48",x"7e",x"bf",x"cd"),
   167 => (x"03",x"a8",x"b7",x"c7"),
   168 => (x"6e",x"87",x"cb",x"c0"),
   169 => (x"c2",x"80",x"c1",x"48"),
   170 => (x"c0",x"58",x"d1",x"f4"),
   171 => (x"4c",x"fe",x"87",x"c2"),
   172 => (x"fd",x"c3",x"4d",x"c1"),
   173 => (x"f8",x"df",x"ff",x"49"),
   174 => (x"c2",x"49",x"70",x"87"),
   175 => (x"87",x"d5",x"02",x"99"),
   176 => (x"bf",x"cd",x"f4",x"c2"),
   177 => (x"87",x"c9",x"c0",x"02"),
   178 => (x"48",x"cd",x"f4",x"c2"),
   179 => (x"c2",x"c0",x"78",x"c0"),
   180 => (x"c1",x"4c",x"fd",x"87"),
   181 => (x"49",x"fa",x"c3",x"4d"),
   182 => (x"87",x"d5",x"df",x"ff"),
   183 => (x"99",x"c2",x"49",x"70"),
   184 => (x"87",x"d9",x"c0",x"02"),
   185 => (x"bf",x"cd",x"f4",x"c2"),
   186 => (x"a8",x"b7",x"c7",x"48"),
   187 => (x"87",x"c9",x"c0",x"03"),
   188 => (x"48",x"cd",x"f4",x"c2"),
   189 => (x"c2",x"c0",x"78",x"c7"),
   190 => (x"c1",x"4c",x"fc",x"87"),
   191 => (x"ac",x"b7",x"c0",x"4d"),
   192 => (x"87",x"d3",x"c0",x"03"),
   193 => (x"c1",x"48",x"66",x"c4"),
   194 => (x"7e",x"70",x"80",x"d8"),
   195 => (x"c0",x"02",x"bf",x"6e"),
   196 => (x"74",x"4b",x"87",x"c5"),
   197 => (x"c0",x"0f",x"73",x"49"),
   198 => (x"1e",x"f0",x"c3",x"1e"),
   199 => (x"f7",x"49",x"da",x"c1"),
   200 => (x"86",x"c8",x"87",x"cb"),
   201 => (x"c0",x"02",x"98",x"70"),
   202 => (x"f4",x"c2",x"87",x"d8"),
   203 => (x"6e",x"7e",x"bf",x"cd"),
   204 => (x"c4",x"91",x"cb",x"49"),
   205 => (x"82",x"71",x"4a",x"66"),
   206 => (x"c5",x"c0",x"02",x"6a"),
   207 => (x"49",x"6e",x"4b",x"87"),
   208 => (x"9d",x"75",x"0f",x"73"),
   209 => (x"87",x"c8",x"c0",x"02"),
   210 => (x"bf",x"cd",x"f4",x"c2"),
   211 => (x"87",x"e1",x"f2",x"49"),
   212 => (x"bf",x"d7",x"cf",x"c2"),
   213 => (x"87",x"dd",x"c0",x"02"),
   214 => (x"87",x"cb",x"c2",x"49"),
   215 => (x"c0",x"02",x"98",x"70"),
   216 => (x"f4",x"c2",x"87",x"d3"),
   217 => (x"f2",x"49",x"bf",x"cd"),
   218 => (x"49",x"c0",x"87",x"c7"),
   219 => (x"c2",x"87",x"e7",x"f3"),
   220 => (x"c0",x"48",x"d7",x"cf"),
   221 => (x"f3",x"8e",x"f8",x"78"),
   222 => (x"5e",x"0e",x"87",x"c1"),
   223 => (x"0e",x"5d",x"5c",x"5b"),
   224 => (x"c2",x"4c",x"71",x"1e"),
   225 => (x"49",x"bf",x"c9",x"f4"),
   226 => (x"4d",x"a1",x"cd",x"c1"),
   227 => (x"69",x"81",x"d1",x"c1"),
   228 => (x"02",x"9c",x"74",x"7e"),
   229 => (x"a5",x"c4",x"87",x"cf"),
   230 => (x"c2",x"7b",x"74",x"4b"),
   231 => (x"49",x"bf",x"c9",x"f4"),
   232 => (x"6e",x"87",x"e0",x"f2"),
   233 => (x"05",x"9c",x"74",x"7b"),
   234 => (x"4b",x"c0",x"87",x"c4"),
   235 => (x"4b",x"c1",x"87",x"c2"),
   236 => (x"e1",x"f2",x"49",x"73"),
   237 => (x"02",x"66",x"d4",x"87"),
   238 => (x"de",x"49",x"87",x"c7"),
   239 => (x"c2",x"4a",x"70",x"87"),
   240 => (x"c2",x"4a",x"c0",x"87"),
   241 => (x"26",x"5a",x"db",x"cf"),
   242 => (x"00",x"87",x"f0",x"f1"),
   243 => (x"00",x"00",x"00",x"00"),
   244 => (x"00",x"00",x"00",x"00"),
   245 => (x"00",x"00",x"00",x"00"),
   246 => (x"1e",x"00",x"00",x"00"),
   247 => (x"c8",x"ff",x"4a",x"71"),
   248 => (x"a1",x"72",x"49",x"bf"),
   249 => (x"1e",x"4f",x"26",x"48"),
   250 => (x"89",x"bf",x"c8",x"ff"),
   251 => (x"c0",x"c0",x"c0",x"fe"),
   252 => (x"01",x"a9",x"c0",x"c0"),
   253 => (x"4a",x"c0",x"87",x"c4"),
   254 => (x"4a",x"c1",x"87",x"c2"),
   255 => (x"4f",x"26",x"48",x"72"),
   256 => (x"dc",x"d3",x"ff",x"1e"),
   257 => (x"49",x"66",x"c4",x"87"),
   258 => (x"02",x"99",x"c0",x"c2"),
   259 => (x"e0",x"c3",x"87",x"cd"),
   260 => (x"de",x"f3",x"c2",x"1e"),
   261 => (x"eb",x"d4",x"ff",x"49"),
   262 => (x"c4",x"86",x"c4",x"87"),
   263 => (x"c0",x"c4",x"49",x"66"),
   264 => (x"87",x"cd",x"02",x"99"),
   265 => (x"c2",x"1e",x"f0",x"c3"),
   266 => (x"ff",x"49",x"de",x"f3"),
   267 => (x"c4",x"87",x"d5",x"d4"),
   268 => (x"49",x"66",x"c4",x"86"),
   269 => (x"71",x"99",x"ff",x"c1"),
   270 => (x"de",x"f3",x"c2",x"1e"),
   271 => (x"c3",x"d4",x"ff",x"49"),
   272 => (x"d4",x"d2",x"ff",x"87"),
   273 => (x"4f",x"26",x"26",x"87"),
   274 => (x"5c",x"5b",x"5e",x"0e"),
   275 => (x"dc",x"ff",x"0e",x"5d"),
   276 => (x"c2",x"7e",x"c0",x"86"),
   277 => (x"49",x"bf",x"d5",x"f4"),
   278 => (x"1e",x"71",x"81",x"c2"),
   279 => (x"4a",x"c6",x"1e",x"72"),
   280 => (x"87",x"c7",x"f2",x"fd"),
   281 => (x"4a",x"26",x"48",x"71"),
   282 => (x"a6",x"c8",x"49",x"26"),
   283 => (x"d5",x"f4",x"c2",x"58"),
   284 => (x"81",x"c4",x"49",x"bf"),
   285 => (x"1e",x"72",x"1e",x"71"),
   286 => (x"f1",x"fd",x"4a",x"c6"),
   287 => (x"48",x"71",x"87",x"ed"),
   288 => (x"49",x"26",x"4a",x"26"),
   289 => (x"c2",x"58",x"a6",x"cc"),
   290 => (x"49",x"bf",x"ee",x"dc"),
   291 => (x"70",x"87",x"d8",x"fd"),
   292 => (x"ce",x"ca",x"02",x"98"),
   293 => (x"49",x"e0",x"c0",x"87"),
   294 => (x"70",x"87",x"c0",x"fd"),
   295 => (x"f2",x"dc",x"c2",x"49"),
   296 => (x"74",x"4c",x"c0",x"59"),
   297 => (x"fe",x"91",x"c4",x"49"),
   298 => (x"4a",x"69",x"81",x"d0"),
   299 => (x"f4",x"c2",x"49",x"74"),
   300 => (x"c4",x"81",x"bf",x"d5"),
   301 => (x"e5",x"f4",x"c2",x"91"),
   302 => (x"9a",x"79",x"72",x"81"),
   303 => (x"72",x"87",x"d2",x"02"),
   304 => (x"71",x"89",x"c1",x"49"),
   305 => (x"c1",x"48",x"6e",x"9a"),
   306 => (x"72",x"7e",x"70",x"80"),
   307 => (x"ee",x"ff",x"05",x"9a"),
   308 => (x"c2",x"84",x"c1",x"87"),
   309 => (x"ff",x"04",x"ac",x"b7"),
   310 => (x"48",x"6e",x"87",x"c9"),
   311 => (x"a8",x"b7",x"fc",x"c0"),
   312 => (x"87",x"ff",x"c8",x"04"),
   313 => (x"4a",x"74",x"4c",x"c0"),
   314 => (x"c4",x"82",x"66",x"c4"),
   315 => (x"e5",x"f4",x"c2",x"92"),
   316 => (x"c8",x"49",x"74",x"82"),
   317 => (x"91",x"c4",x"81",x"66"),
   318 => (x"81",x"e5",x"f4",x"c2"),
   319 => (x"49",x"69",x"4a",x"6a"),
   320 => (x"4b",x"74",x"b9",x"72"),
   321 => (x"bf",x"d5",x"f4",x"c2"),
   322 => (x"c2",x"93",x"c4",x"83"),
   323 => (x"6b",x"83",x"e5",x"f4"),
   324 => (x"71",x"48",x"72",x"ba"),
   325 => (x"58",x"a6",x"d0",x"98"),
   326 => (x"f4",x"c2",x"49",x"74"),
   327 => (x"c4",x"81",x"bf",x"d5"),
   328 => (x"e5",x"f4",x"c2",x"91"),
   329 => (x"d0",x"7e",x"69",x"81"),
   330 => (x"78",x"c0",x"48",x"a6"),
   331 => (x"df",x"49",x"66",x"cc"),
   332 => (x"c0",x"c7",x"02",x"29"),
   333 => (x"c0",x"4a",x"74",x"87"),
   334 => (x"66",x"d0",x"92",x"e0"),
   335 => (x"48",x"ff",x"c0",x"82"),
   336 => (x"4a",x"70",x"88",x"72"),
   337 => (x"c0",x"48",x"a6",x"d4"),
   338 => (x"c0",x"80",x"c4",x"78"),
   339 => (x"df",x"49",x"6e",x"78"),
   340 => (x"a6",x"e0",x"c0",x"29"),
   341 => (x"d1",x"f4",x"c2",x"59"),
   342 => (x"72",x"78",x"c1",x"48"),
   343 => (x"b7",x"31",x"c3",x"49"),
   344 => (x"c0",x"b1",x"72",x"2a"),
   345 => (x"91",x"c4",x"99",x"ff"),
   346 => (x"4d",x"c5",x"de",x"c2"),
   347 => (x"4b",x"6d",x"85",x"71"),
   348 => (x"c0",x"c0",x"c4",x"49"),
   349 => (x"f3",x"c0",x"02",x"99"),
   350 => (x"02",x"66",x"dc",x"87"),
   351 => (x"80",x"c8",x"87",x"c8"),
   352 => (x"c5",x"78",x"40",x"c0"),
   353 => (x"f4",x"c2",x"87",x"ef"),
   354 => (x"78",x"c1",x"48",x"d9"),
   355 => (x"bf",x"dd",x"f4",x"c2"),
   356 => (x"87",x"e1",x"c5",x"05"),
   357 => (x"f8",x"1e",x"d8",x"c1"),
   358 => (x"e3",x"f9",x"49",x"a0"),
   359 => (x"1e",x"d8",x"c5",x"87"),
   360 => (x"49",x"d1",x"f4",x"c2"),
   361 => (x"c8",x"87",x"d9",x"f9"),
   362 => (x"87",x"c9",x"c5",x"86"),
   363 => (x"d8",x"02",x"66",x"dc"),
   364 => (x"c2",x"49",x"73",x"87"),
   365 => (x"02",x"99",x"c0",x"c0"),
   366 => (x"d0",x"87",x"c3",x"c0"),
   367 => (x"48",x"6d",x"2b",x"b7"),
   368 => (x"98",x"ff",x"ff",x"fd"),
   369 => (x"fa",x"c0",x"7d",x"70"),
   370 => (x"d9",x"f4",x"c2",x"87"),
   371 => (x"f2",x"c0",x"02",x"bf"),
   372 => (x"d0",x"48",x"73",x"87"),
   373 => (x"e4",x"c0",x"28",x"b7"),
   374 => (x"98",x"70",x"58",x"a6"),
   375 => (x"87",x"e3",x"c0",x"02"),
   376 => (x"bf",x"e1",x"f4",x"c2"),
   377 => (x"c0",x"e0",x"c0",x"49"),
   378 => (x"ca",x"c0",x"02",x"99"),
   379 => (x"c0",x"49",x"70",x"87"),
   380 => (x"02",x"99",x"c0",x"e0"),
   381 => (x"6d",x"87",x"cc",x"c0"),
   382 => (x"c0",x"c0",x"c2",x"48"),
   383 => (x"c0",x"7d",x"70",x"b0"),
   384 => (x"73",x"4b",x"66",x"e0"),
   385 => (x"c0",x"c0",x"c8",x"49"),
   386 => (x"c7",x"c2",x"02",x"99"),
   387 => (x"e1",x"f4",x"c2",x"87"),
   388 => (x"c0",x"cc",x"4a",x"bf"),
   389 => (x"cf",x"c0",x"02",x"9a"),
   390 => (x"8a",x"c0",x"c4",x"87"),
   391 => (x"87",x"d8",x"c0",x"02"),
   392 => (x"f9",x"c0",x"02",x"8a"),
   393 => (x"87",x"dd",x"c1",x"87"),
   394 => (x"ff",x"c3",x"49",x"73"),
   395 => (x"c2",x"91",x"c2",x"99"),
   396 => (x"11",x"81",x"f9",x"dd"),
   397 => (x"87",x"dc",x"c1",x"4b"),
   398 => (x"ff",x"c3",x"49",x"73"),
   399 => (x"c2",x"91",x"c2",x"99"),
   400 => (x"c1",x"81",x"f9",x"dd"),
   401 => (x"dc",x"4b",x"11",x"81"),
   402 => (x"c8",x"c0",x"02",x"66"),
   403 => (x"48",x"a6",x"d8",x"87"),
   404 => (x"ff",x"c0",x"78",x"d2"),
   405 => (x"48",x"a6",x"d4",x"87"),
   406 => (x"c0",x"78",x"d2",x"c4"),
   407 => (x"49",x"73",x"87",x"f6"),
   408 => (x"c2",x"99",x"ff",x"c3"),
   409 => (x"f9",x"dd",x"c2",x"91"),
   410 => (x"11",x"81",x"c1",x"81"),
   411 => (x"02",x"66",x"dc",x"4b"),
   412 => (x"d8",x"87",x"c9",x"c0"),
   413 => (x"d9",x"c1",x"48",x"a6"),
   414 => (x"87",x"d8",x"c0",x"78"),
   415 => (x"c5",x"48",x"a6",x"d4"),
   416 => (x"cf",x"c0",x"78",x"d9"),
   417 => (x"c3",x"49",x"73",x"87"),
   418 => (x"91",x"c2",x"99",x"ff"),
   419 => (x"81",x"f9",x"dd",x"c2"),
   420 => (x"4b",x"11",x"81",x"c1"),
   421 => (x"c0",x"02",x"66",x"dc"),
   422 => (x"49",x"73",x"87",x"dc"),
   423 => (x"fc",x"c7",x"b9",x"ff"),
   424 => (x"48",x"71",x"99",x"c0"),
   425 => (x"bf",x"e1",x"f4",x"c2"),
   426 => (x"e5",x"f4",x"c2",x"98"),
   427 => (x"9b",x"ff",x"c3",x"58"),
   428 => (x"c0",x"b3",x"c0",x"c4"),
   429 => (x"49",x"73",x"87",x"d4"),
   430 => (x"99",x"c0",x"fc",x"c7"),
   431 => (x"f4",x"c2",x"48",x"71"),
   432 => (x"c2",x"b0",x"bf",x"e1"),
   433 => (x"c3",x"58",x"e5",x"f4"),
   434 => (x"66",x"d4",x"9b",x"ff"),
   435 => (x"87",x"ca",x"c0",x"02"),
   436 => (x"d1",x"f4",x"c2",x"1e"),
   437 => (x"87",x"e8",x"f4",x"49"),
   438 => (x"1e",x"73",x"86",x"c4"),
   439 => (x"49",x"d1",x"f4",x"c2"),
   440 => (x"c4",x"87",x"dd",x"f4"),
   441 => (x"02",x"66",x"d8",x"86"),
   442 => (x"1e",x"87",x"ca",x"c0"),
   443 => (x"49",x"d1",x"f4",x"c2"),
   444 => (x"c4",x"87",x"cd",x"f4"),
   445 => (x"48",x"66",x"cc",x"86"),
   446 => (x"a6",x"d0",x"30",x"c1"),
   447 => (x"c1",x"48",x"6e",x"58"),
   448 => (x"d0",x"7e",x"70",x"30"),
   449 => (x"80",x"c1",x"48",x"66"),
   450 => (x"c0",x"58",x"a6",x"d4"),
   451 => (x"04",x"a8",x"b7",x"e0"),
   452 => (x"c1",x"87",x"d9",x"f8"),
   453 => (x"ac",x"b7",x"c2",x"84"),
   454 => (x"87",x"ca",x"f7",x"04"),
   455 => (x"48",x"d5",x"f4",x"c2"),
   456 => (x"ff",x"78",x"66",x"c4"),
   457 => (x"4d",x"26",x"8e",x"dc"),
   458 => (x"4b",x"26",x"4c",x"26"),
   459 => (x"00",x"00",x"4f",x"26"),
   460 => (x"c0",x"1e",x"00",x"00"),
   461 => (x"c4",x"49",x"72",x"4a"),
   462 => (x"e5",x"f4",x"c2",x"91"),
   463 => (x"c1",x"79",x"ff",x"81"),
   464 => (x"aa",x"b7",x"c6",x"82"),
   465 => (x"c2",x"87",x"ee",x"04"),
   466 => (x"c0",x"48",x"d5",x"f4"),
   467 => (x"80",x"c8",x"78",x"40"),
   468 => (x"4f",x"26",x"78",x"c0"),
   469 => (x"71",x"1e",x"73",x"1e"),
   470 => (x"f5",x"dd",x"c2",x"4b"),
   471 => (x"87",x"c9",x"05",x"bf"),
   472 => (x"48",x"f5",x"dd",x"c2"),
   473 => (x"c9",x"ff",x"78",x"c1"),
   474 => (x"87",x"dc",x"f3",x"87"),
   475 => (x"c8",x"ff",x"49",x"73"),
   476 => (x"f5",x"fe",x"87",x"fc"),
   477 => (x"00",x"00",x"00",x"87"),
   478 => (x"f2",x"eb",x"f4",x"00"),
   479 => (x"04",x"06",x"05",x"f5"),
   480 => (x"83",x"0b",x"03",x"0c"),
   481 => (x"fc",x"00",x"66",x"0a"),
   482 => (x"da",x"00",x"5a",x"00"),
   483 => (x"94",x"80",x"00",x"00"),
   484 => (x"78",x"80",x"05",x"08"),
   485 => (x"01",x"80",x"02",x"00"),
   486 => (x"09",x"80",x"03",x"00"),
   487 => (x"00",x"80",x"04",x"00"),
   488 => (x"91",x"80",x"01",x"00"),
   489 => (x"04",x"00",x"26",x"08"),
   490 => (x"00",x"00",x"1d",x"00"),
   491 => (x"00",x"00",x"1c",x"00"),
   492 => (x"0c",x"00",x"25",x"00"),
   493 => (x"00",x"00",x"1a",x"00"),
   494 => (x"00",x"00",x"1b",x"00"),
   495 => (x"00",x"00",x"24",x"00"),
   496 => (x"00",x"01",x"12",x"00"),
   497 => (x"03",x"00",x"2e",x"00"),
   498 => (x"00",x"00",x"2d",x"00"),
   499 => (x"00",x"00",x"23",x"00"),
   500 => (x"0b",x"00",x"36",x"00"),
   501 => (x"00",x"00",x"21",x"00"),
   502 => (x"00",x"00",x"2b",x"00"),
   503 => (x"00",x"00",x"2c",x"00"),
   504 => (x"00",x"00",x"22",x"00"),
   505 => (x"6c",x"00",x"3d",x"00"),
   506 => (x"00",x"00",x"35",x"00"),
   507 => (x"00",x"00",x"34",x"00"),
   508 => (x"75",x"00",x"3e",x"00"),
   509 => (x"00",x"00",x"32",x"00"),
   510 => (x"00",x"00",x"33",x"00"),
   511 => (x"6b",x"00",x"3c",x"00"),
   512 => (x"00",x"00",x"2a",x"00"),
   513 => (x"01",x"00",x"46",x"00"),
   514 => (x"73",x"00",x"43",x"00"),
   515 => (x"69",x"00",x"3b",x"00"),
   516 => (x"09",x"00",x"45",x"00"),
   517 => (x"70",x"00",x"3a",x"00"),
   518 => (x"72",x"00",x"42",x"00"),
   519 => (x"74",x"00",x"44",x"00"),
   520 => (x"00",x"00",x"31",x"00"),
   521 => (x"00",x"00",x"55",x"00"),
   522 => (x"7c",x"00",x"4d",x"00"),
   523 => (x"7a",x"00",x"4b",x"00"),
   524 => (x"00",x"00",x"7b",x"00"),
   525 => (x"71",x"00",x"49",x"00"),
   526 => (x"84",x"00",x"4c",x"00"),
   527 => (x"77",x"00",x"54",x"00"),
   528 => (x"00",x"00",x"41",x"00"),
   529 => (x"00",x"00",x"61",x"00"),
   530 => (x"7c",x"00",x"5b",x"00"),
   531 => (x"00",x"00",x"52",x"00"),
   532 => (x"00",x"00",x"f1",x"00"),
   533 => (x"00",x"02",x"59",x"00"),
   534 => (x"5d",x"00",x"0e",x"00"),
   535 => (x"00",x"00",x"5d",x"00"),
   536 => (x"79",x"00",x"4a",x"00"),
   537 => (x"05",x"00",x"16",x"00"),
   538 => (x"07",x"00",x"76",x"00"),
   539 => (x"0d",x"00",x"0d",x"00"),
   540 => (x"06",x"00",x"1e",x"00"),
   541 => (x"00",x"00",x"29",x"00"),
   542 => (x"00",x"04",x"14",x"00"),
   543 => (x"00",x"00",x"15",x"00"),
   544 => (x"00",x"40",x"00",x"00"),
   545 => (x"00",x"40",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

