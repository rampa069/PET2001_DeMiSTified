
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"f5",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"d8",x"f5",x"c2"),
    14 => (x"48",x"c8",x"e2",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"db",x"df"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"9a",x"72",x"1e",x"73"),
    47 => (x"87",x"e7",x"c0",x"02"),
    48 => (x"4b",x"c1",x"48",x"c0"),
    49 => (x"d1",x"06",x"a9",x"72"),
    50 => (x"06",x"82",x"72",x"87"),
    51 => (x"83",x"73",x"87",x"c9"),
    52 => (x"f4",x"01",x"a9",x"72"),
    53 => (x"c1",x"87",x"c3",x"87"),
    54 => (x"a9",x"72",x"3a",x"b2"),
    55 => (x"80",x"73",x"89",x"03"),
    56 => (x"2b",x"2a",x"c1",x"07"),
    57 => (x"26",x"87",x"f3",x"05"),
    58 => (x"1e",x"4f",x"26",x"4b"),
    59 => (x"4d",x"c4",x"1e",x"75"),
    60 => (x"04",x"a1",x"b7",x"71"),
    61 => (x"81",x"c1",x"b9",x"ff"),
    62 => (x"72",x"07",x"bd",x"c3"),
    63 => (x"ff",x"04",x"a2",x"b7"),
    64 => (x"c1",x"82",x"c1",x"ba"),
    65 => (x"ee",x"fe",x"07",x"bd"),
    66 => (x"04",x"2d",x"c1",x"87"),
    67 => (x"80",x"c1",x"b8",x"ff"),
    68 => (x"ff",x"04",x"2d",x"07"),
    69 => (x"07",x"81",x"c1",x"b9"),
    70 => (x"4f",x"26",x"4d",x"26"),
    71 => (x"c4",x"4a",x"71",x"1e"),
    72 => (x"c1",x"48",x"49",x"66"),
    73 => (x"58",x"a6",x"c8",x"88"),
    74 => (x"d6",x"02",x"99",x"71"),
    75 => (x"48",x"d4",x"ff",x"87"),
    76 => (x"68",x"78",x"ff",x"c3"),
    77 => (x"49",x"66",x"c4",x"52"),
    78 => (x"c8",x"88",x"c1",x"48"),
    79 => (x"99",x"71",x"58",x"a6"),
    80 => (x"26",x"87",x"ea",x"05"),
    81 => (x"1e",x"73",x"1e",x"4f"),
    82 => (x"c3",x"4b",x"d4",x"ff"),
    83 => (x"4a",x"6b",x"7b",x"ff"),
    84 => (x"6b",x"7b",x"ff",x"c3"),
    85 => (x"72",x"32",x"c8",x"49"),
    86 => (x"7b",x"ff",x"c3",x"b1"),
    87 => (x"31",x"c8",x"4a",x"6b"),
    88 => (x"ff",x"c3",x"b2",x"71"),
    89 => (x"c8",x"49",x"6b",x"7b"),
    90 => (x"71",x"b1",x"72",x"32"),
    91 => (x"26",x"87",x"c4",x"48"),
    92 => (x"26",x"4c",x"26",x"4d"),
    93 => (x"0e",x"4f",x"26",x"4b"),
    94 => (x"5d",x"5c",x"5b",x"5e"),
    95 => (x"ff",x"4a",x"71",x"0e"),
    96 => (x"49",x"72",x"4c",x"d4"),
    97 => (x"71",x"99",x"ff",x"c3"),
    98 => (x"c8",x"e2",x"c2",x"7c"),
    99 => (x"87",x"c8",x"05",x"bf"),
   100 => (x"c9",x"48",x"66",x"d0"),
   101 => (x"58",x"a6",x"d4",x"30"),
   102 => (x"d8",x"49",x"66",x"d0"),
   103 => (x"99",x"ff",x"c3",x"29"),
   104 => (x"66",x"d0",x"7c",x"71"),
   105 => (x"c3",x"29",x"d0",x"49"),
   106 => (x"7c",x"71",x"99",x"ff"),
   107 => (x"c8",x"49",x"66",x"d0"),
   108 => (x"99",x"ff",x"c3",x"29"),
   109 => (x"66",x"d0",x"7c",x"71"),
   110 => (x"99",x"ff",x"c3",x"49"),
   111 => (x"49",x"72",x"7c",x"71"),
   112 => (x"ff",x"c3",x"29",x"d0"),
   113 => (x"6c",x"7c",x"71",x"99"),
   114 => (x"ff",x"f0",x"c9",x"4b"),
   115 => (x"ab",x"ff",x"c3",x"4d"),
   116 => (x"c3",x"87",x"d0",x"05"),
   117 => (x"4b",x"6c",x"7c",x"ff"),
   118 => (x"c6",x"02",x"8d",x"c1"),
   119 => (x"ab",x"ff",x"c3",x"87"),
   120 => (x"73",x"87",x"f0",x"02"),
   121 => (x"87",x"c7",x"fe",x"48"),
   122 => (x"ff",x"49",x"c0",x"1e"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"c3",x"81",x"c1",x"78"),
   125 => (x"04",x"a9",x"b7",x"c8"),
   126 => (x"4f",x"26",x"87",x"f1"),
   127 => (x"e7",x"1e",x"73",x"1e"),
   128 => (x"df",x"f8",x"c4",x"87"),
   129 => (x"c0",x"1e",x"c0",x"4b"),
   130 => (x"f7",x"c1",x"f0",x"ff"),
   131 => (x"87",x"e7",x"fd",x"49"),
   132 => (x"a8",x"c1",x"86",x"c4"),
   133 => (x"87",x"ea",x"c0",x"05"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"c0",x"c1",x"78",x"ff"),
   136 => (x"c0",x"c0",x"c0",x"c0"),
   137 => (x"f0",x"e1",x"c0",x"1e"),
   138 => (x"fd",x"49",x"e9",x"c1"),
   139 => (x"86",x"c4",x"87",x"c9"),
   140 => (x"ca",x"05",x"98",x"70"),
   141 => (x"48",x"d4",x"ff",x"87"),
   142 => (x"c1",x"78",x"ff",x"c3"),
   143 => (x"fe",x"87",x"cb",x"48"),
   144 => (x"8b",x"c1",x"87",x"e6"),
   145 => (x"87",x"fd",x"fe",x"05"),
   146 => (x"e6",x"fc",x"48",x"c0"),
   147 => (x"1e",x"73",x"1e",x"87"),
   148 => (x"c3",x"48",x"d4",x"ff"),
   149 => (x"4b",x"d3",x"78",x"ff"),
   150 => (x"ff",x"c0",x"1e",x"c0"),
   151 => (x"49",x"c1",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d4",x"fc"),
   153 => (x"05",x"98",x"70",x"86"),
   154 => (x"d4",x"ff",x"87",x"ca"),
   155 => (x"78",x"ff",x"c3",x"48"),
   156 => (x"87",x"cb",x"48",x"c1"),
   157 => (x"c1",x"87",x"f1",x"fd"),
   158 => (x"db",x"ff",x"05",x"8b"),
   159 => (x"fb",x"48",x"c0",x"87"),
   160 => (x"5e",x"0e",x"87",x"f1"),
   161 => (x"ff",x"0e",x"5c",x"5b"),
   162 => (x"db",x"fd",x"4c",x"d4"),
   163 => (x"1e",x"ea",x"c6",x"87"),
   164 => (x"c1",x"f0",x"e1",x"c0"),
   165 => (x"de",x"fb",x"49",x"c8"),
   166 => (x"c1",x"86",x"c4",x"87"),
   167 => (x"87",x"c8",x"02",x"a8"),
   168 => (x"c0",x"87",x"ea",x"fe"),
   169 => (x"87",x"e2",x"c1",x"48"),
   170 => (x"70",x"87",x"da",x"fa"),
   171 => (x"ff",x"ff",x"cf",x"49"),
   172 => (x"a9",x"ea",x"c6",x"99"),
   173 => (x"fe",x"87",x"c8",x"02"),
   174 => (x"48",x"c0",x"87",x"d3"),
   175 => (x"c3",x"87",x"cb",x"c1"),
   176 => (x"f1",x"c0",x"7c",x"ff"),
   177 => (x"87",x"f4",x"fc",x"4b"),
   178 => (x"c0",x"02",x"98",x"70"),
   179 => (x"1e",x"c0",x"87",x"eb"),
   180 => (x"c1",x"f0",x"ff",x"c0"),
   181 => (x"de",x"fa",x"49",x"fa"),
   182 => (x"70",x"86",x"c4",x"87"),
   183 => (x"87",x"d9",x"05",x"98"),
   184 => (x"6c",x"7c",x"ff",x"c3"),
   185 => (x"7c",x"ff",x"c3",x"49"),
   186 => (x"c1",x"7c",x"7c",x"7c"),
   187 => (x"c4",x"02",x"99",x"c0"),
   188 => (x"d5",x"48",x"c1",x"87"),
   189 => (x"d1",x"48",x"c0",x"87"),
   190 => (x"05",x"ab",x"c2",x"87"),
   191 => (x"48",x"c0",x"87",x"c4"),
   192 => (x"8b",x"c1",x"87",x"c8"),
   193 => (x"87",x"fd",x"fe",x"05"),
   194 => (x"e4",x"f9",x"48",x"c0"),
   195 => (x"1e",x"73",x"1e",x"87"),
   196 => (x"48",x"c8",x"e2",x"c2"),
   197 => (x"4b",x"c7",x"78",x"c1"),
   198 => (x"c2",x"48",x"d0",x"ff"),
   199 => (x"87",x"c8",x"fb",x"78"),
   200 => (x"c3",x"48",x"d0",x"ff"),
   201 => (x"c0",x"1e",x"c0",x"78"),
   202 => (x"c0",x"c1",x"d0",x"e5"),
   203 => (x"87",x"c7",x"f9",x"49"),
   204 => (x"a8",x"c1",x"86",x"c4"),
   205 => (x"4b",x"87",x"c1",x"05"),
   206 => (x"c5",x"05",x"ab",x"c2"),
   207 => (x"c0",x"48",x"c0",x"87"),
   208 => (x"8b",x"c1",x"87",x"f9"),
   209 => (x"87",x"d0",x"ff",x"05"),
   210 => (x"c2",x"87",x"f7",x"fc"),
   211 => (x"70",x"58",x"cc",x"e2"),
   212 => (x"87",x"cd",x"05",x"98"),
   213 => (x"ff",x"c0",x"1e",x"c1"),
   214 => (x"49",x"d0",x"c1",x"f0"),
   215 => (x"c4",x"87",x"d8",x"f8"),
   216 => (x"48",x"d4",x"ff",x"86"),
   217 => (x"c2",x"78",x"ff",x"c3"),
   218 => (x"e2",x"c2",x"87",x"fc"),
   219 => (x"d0",x"ff",x"58",x"d0"),
   220 => (x"ff",x"78",x"c2",x"48"),
   221 => (x"ff",x"c3",x"48",x"d4"),
   222 => (x"f7",x"48",x"c1",x"78"),
   223 => (x"5e",x"0e",x"87",x"f5"),
   224 => (x"0e",x"5d",x"5c",x"5b"),
   225 => (x"4c",x"c0",x"4b",x"71"),
   226 => (x"df",x"cd",x"ee",x"c5"),
   227 => (x"48",x"d4",x"ff",x"4a"),
   228 => (x"68",x"78",x"ff",x"c3"),
   229 => (x"a9",x"fe",x"c3",x"49"),
   230 => (x"87",x"fd",x"c0",x"05"),
   231 => (x"9b",x"73",x"4d",x"70"),
   232 => (x"d0",x"87",x"cc",x"02"),
   233 => (x"49",x"73",x"1e",x"66"),
   234 => (x"c4",x"87",x"f1",x"f5"),
   235 => (x"ff",x"87",x"d6",x"86"),
   236 => (x"d1",x"c4",x"48",x"d0"),
   237 => (x"7d",x"ff",x"c3",x"78"),
   238 => (x"c1",x"48",x"66",x"d0"),
   239 => (x"58",x"a6",x"d4",x"88"),
   240 => (x"f0",x"05",x"98",x"70"),
   241 => (x"48",x"d4",x"ff",x"87"),
   242 => (x"78",x"78",x"ff",x"c3"),
   243 => (x"c5",x"05",x"9b",x"73"),
   244 => (x"48",x"d0",x"ff",x"87"),
   245 => (x"4a",x"c1",x"78",x"d0"),
   246 => (x"05",x"8a",x"c1",x"4c"),
   247 => (x"74",x"87",x"ee",x"fe"),
   248 => (x"87",x"cb",x"f6",x"48"),
   249 => (x"71",x"1e",x"73",x"1e"),
   250 => (x"ff",x"4b",x"c0",x"4a"),
   251 => (x"ff",x"c3",x"48",x"d4"),
   252 => (x"48",x"d0",x"ff",x"78"),
   253 => (x"ff",x"78",x"c3",x"c4"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"c0",x"1e",x"72",x"78"),
   256 => (x"d1",x"c1",x"f0",x"ff"),
   257 => (x"87",x"ef",x"f5",x"49"),
   258 => (x"98",x"70",x"86",x"c4"),
   259 => (x"c8",x"87",x"d2",x"05"),
   260 => (x"66",x"cc",x"1e",x"c0"),
   261 => (x"87",x"e6",x"fd",x"49"),
   262 => (x"4b",x"70",x"86",x"c4"),
   263 => (x"c2",x"48",x"d0",x"ff"),
   264 => (x"f5",x"48",x"73",x"78"),
   265 => (x"5e",x"0e",x"87",x"cd"),
   266 => (x"0e",x"5d",x"5c",x"5b"),
   267 => (x"ff",x"c0",x"1e",x"c0"),
   268 => (x"49",x"c9",x"c1",x"f0"),
   269 => (x"d2",x"87",x"c0",x"f5"),
   270 => (x"d0",x"e2",x"c2",x"1e"),
   271 => (x"87",x"fe",x"fc",x"49"),
   272 => (x"4c",x"c0",x"86",x"c8"),
   273 => (x"b7",x"d2",x"84",x"c1"),
   274 => (x"87",x"f8",x"04",x"ac"),
   275 => (x"97",x"d0",x"e2",x"c2"),
   276 => (x"c0",x"c3",x"49",x"bf"),
   277 => (x"a9",x"c0",x"c1",x"99"),
   278 => (x"87",x"e7",x"c0",x"05"),
   279 => (x"97",x"d7",x"e2",x"c2"),
   280 => (x"31",x"d0",x"49",x"bf"),
   281 => (x"97",x"d8",x"e2",x"c2"),
   282 => (x"32",x"c8",x"4a",x"bf"),
   283 => (x"e2",x"c2",x"b1",x"72"),
   284 => (x"4a",x"bf",x"97",x"d9"),
   285 => (x"cf",x"4c",x"71",x"b1"),
   286 => (x"9c",x"ff",x"ff",x"ff"),
   287 => (x"34",x"ca",x"84",x"c1"),
   288 => (x"c2",x"87",x"e7",x"c1"),
   289 => (x"bf",x"97",x"d9",x"e2"),
   290 => (x"c6",x"31",x"c1",x"49"),
   291 => (x"da",x"e2",x"c2",x"99"),
   292 => (x"c7",x"4a",x"bf",x"97"),
   293 => (x"b1",x"72",x"2a",x"b7"),
   294 => (x"97",x"d5",x"e2",x"c2"),
   295 => (x"cf",x"4d",x"4a",x"bf"),
   296 => (x"d6",x"e2",x"c2",x"9d"),
   297 => (x"c3",x"4a",x"bf",x"97"),
   298 => (x"c2",x"32",x"ca",x"9a"),
   299 => (x"bf",x"97",x"d7",x"e2"),
   300 => (x"73",x"33",x"c2",x"4b"),
   301 => (x"d8",x"e2",x"c2",x"b2"),
   302 => (x"c3",x"4b",x"bf",x"97"),
   303 => (x"b7",x"c6",x"9b",x"c0"),
   304 => (x"c2",x"b2",x"73",x"2b"),
   305 => (x"71",x"48",x"c1",x"81"),
   306 => (x"c1",x"49",x"70",x"30"),
   307 => (x"70",x"30",x"75",x"48"),
   308 => (x"c1",x"4c",x"72",x"4d"),
   309 => (x"c8",x"94",x"71",x"84"),
   310 => (x"06",x"ad",x"b7",x"c0"),
   311 => (x"34",x"c1",x"87",x"cc"),
   312 => (x"c0",x"c8",x"2d",x"b7"),
   313 => (x"ff",x"01",x"ad",x"b7"),
   314 => (x"48",x"74",x"87",x"f4"),
   315 => (x"0e",x"87",x"c0",x"f2"),
   316 => (x"5d",x"5c",x"5b",x"5e"),
   317 => (x"c2",x"86",x"f8",x"0e"),
   318 => (x"c0",x"48",x"f6",x"ea"),
   319 => (x"ee",x"e2",x"c2",x"78"),
   320 => (x"fb",x"49",x"c0",x"1e"),
   321 => (x"86",x"c4",x"87",x"de"),
   322 => (x"c5",x"05",x"98",x"70"),
   323 => (x"c9",x"48",x"c0",x"87"),
   324 => (x"4d",x"c0",x"87",x"ce"),
   325 => (x"ef",x"c0",x"7e",x"c1"),
   326 => (x"c2",x"49",x"bf",x"d8"),
   327 => (x"71",x"4a",x"e4",x"e3"),
   328 => (x"c4",x"ed",x"4b",x"c8"),
   329 => (x"05",x"98",x"70",x"87"),
   330 => (x"7e",x"c0",x"87",x"c2"),
   331 => (x"bf",x"d4",x"ef",x"c0"),
   332 => (x"c0",x"e4",x"c2",x"49"),
   333 => (x"4b",x"c8",x"71",x"4a"),
   334 => (x"70",x"87",x"ee",x"ec"),
   335 => (x"87",x"c2",x"05",x"98"),
   336 => (x"02",x"6e",x"7e",x"c0"),
   337 => (x"c2",x"87",x"fd",x"c0"),
   338 => (x"4d",x"bf",x"f4",x"e9"),
   339 => (x"9f",x"ec",x"ea",x"c2"),
   340 => (x"c5",x"48",x"7e",x"bf"),
   341 => (x"05",x"a8",x"ea",x"d6"),
   342 => (x"e9",x"c2",x"87",x"c7"),
   343 => (x"ce",x"4d",x"bf",x"f4"),
   344 => (x"ca",x"48",x"6e",x"87"),
   345 => (x"02",x"a8",x"d5",x"e9"),
   346 => (x"48",x"c0",x"87",x"c5"),
   347 => (x"c2",x"87",x"f1",x"c7"),
   348 => (x"75",x"1e",x"ee",x"e2"),
   349 => (x"87",x"ec",x"f9",x"49"),
   350 => (x"98",x"70",x"86",x"c4"),
   351 => (x"c0",x"87",x"c5",x"05"),
   352 => (x"87",x"dc",x"c7",x"48"),
   353 => (x"bf",x"d4",x"ef",x"c0"),
   354 => (x"c0",x"e4",x"c2",x"49"),
   355 => (x"4b",x"c8",x"71",x"4a"),
   356 => (x"70",x"87",x"d6",x"eb"),
   357 => (x"87",x"c8",x"05",x"98"),
   358 => (x"48",x"f6",x"ea",x"c2"),
   359 => (x"87",x"da",x"78",x"c1"),
   360 => (x"bf",x"d8",x"ef",x"c0"),
   361 => (x"e4",x"e3",x"c2",x"49"),
   362 => (x"4b",x"c8",x"71",x"4a"),
   363 => (x"70",x"87",x"fa",x"ea"),
   364 => (x"c5",x"c0",x"02",x"98"),
   365 => (x"c6",x"48",x"c0",x"87"),
   366 => (x"ea",x"c2",x"87",x"e6"),
   367 => (x"49",x"bf",x"97",x"ec"),
   368 => (x"05",x"a9",x"d5",x"c1"),
   369 => (x"c2",x"87",x"cd",x"c0"),
   370 => (x"bf",x"97",x"ed",x"ea"),
   371 => (x"a9",x"ea",x"c2",x"49"),
   372 => (x"87",x"c5",x"c0",x"02"),
   373 => (x"c7",x"c6",x"48",x"c0"),
   374 => (x"ee",x"e2",x"c2",x"87"),
   375 => (x"48",x"7e",x"bf",x"97"),
   376 => (x"02",x"a8",x"e9",x"c3"),
   377 => (x"6e",x"87",x"ce",x"c0"),
   378 => (x"a8",x"eb",x"c3",x"48"),
   379 => (x"87",x"c5",x"c0",x"02"),
   380 => (x"eb",x"c5",x"48",x"c0"),
   381 => (x"f9",x"e2",x"c2",x"87"),
   382 => (x"99",x"49",x"bf",x"97"),
   383 => (x"87",x"cc",x"c0",x"05"),
   384 => (x"97",x"fa",x"e2",x"c2"),
   385 => (x"a9",x"c2",x"49",x"bf"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"cf",x"c5",x"48",x"c0"),
   388 => (x"fb",x"e2",x"c2",x"87"),
   389 => (x"c2",x"48",x"bf",x"97"),
   390 => (x"70",x"58",x"f2",x"ea"),
   391 => (x"88",x"c1",x"48",x"4c"),
   392 => (x"58",x"f6",x"ea",x"c2"),
   393 => (x"97",x"fc",x"e2",x"c2"),
   394 => (x"81",x"75",x"49",x"bf"),
   395 => (x"97",x"fd",x"e2",x"c2"),
   396 => (x"32",x"c8",x"4a",x"bf"),
   397 => (x"c2",x"7e",x"a1",x"72"),
   398 => (x"6e",x"48",x"c3",x"ef"),
   399 => (x"fe",x"e2",x"c2",x"78"),
   400 => (x"c8",x"48",x"bf",x"97"),
   401 => (x"ea",x"c2",x"58",x"a6"),
   402 => (x"c2",x"02",x"bf",x"f6"),
   403 => (x"ef",x"c0",x"87",x"d4"),
   404 => (x"c2",x"49",x"bf",x"d4"),
   405 => (x"71",x"4a",x"c0",x"e4"),
   406 => (x"cc",x"e8",x"4b",x"c8"),
   407 => (x"02",x"98",x"70",x"87"),
   408 => (x"c0",x"87",x"c5",x"c0"),
   409 => (x"87",x"f8",x"c3",x"48"),
   410 => (x"bf",x"ee",x"ea",x"c2"),
   411 => (x"d7",x"ef",x"c2",x"4c"),
   412 => (x"d3",x"e3",x"c2",x"5c"),
   413 => (x"c8",x"49",x"bf",x"97"),
   414 => (x"d2",x"e3",x"c2",x"31"),
   415 => (x"a1",x"4a",x"bf",x"97"),
   416 => (x"d4",x"e3",x"c2",x"49"),
   417 => (x"d0",x"4a",x"bf",x"97"),
   418 => (x"49",x"a1",x"72",x"32"),
   419 => (x"97",x"d5",x"e3",x"c2"),
   420 => (x"32",x"d8",x"4a",x"bf"),
   421 => (x"c4",x"49",x"a1",x"72"),
   422 => (x"ef",x"c2",x"91",x"66"),
   423 => (x"c2",x"81",x"bf",x"c3"),
   424 => (x"c2",x"59",x"cb",x"ef"),
   425 => (x"bf",x"97",x"db",x"e3"),
   426 => (x"c2",x"32",x"c8",x"4a"),
   427 => (x"bf",x"97",x"da",x"e3"),
   428 => (x"c2",x"4a",x"a2",x"4b"),
   429 => (x"bf",x"97",x"dc",x"e3"),
   430 => (x"73",x"33",x"d0",x"4b"),
   431 => (x"e3",x"c2",x"4a",x"a2"),
   432 => (x"4b",x"bf",x"97",x"dd"),
   433 => (x"33",x"d8",x"9b",x"cf"),
   434 => (x"c2",x"4a",x"a2",x"73"),
   435 => (x"c2",x"5a",x"cf",x"ef"),
   436 => (x"4a",x"bf",x"cb",x"ef"),
   437 => (x"92",x"74",x"8a",x"c2"),
   438 => (x"48",x"cf",x"ef",x"c2"),
   439 => (x"c1",x"78",x"a1",x"72"),
   440 => (x"e3",x"c2",x"87",x"ca"),
   441 => (x"49",x"bf",x"97",x"c0"),
   442 => (x"e2",x"c2",x"31",x"c8"),
   443 => (x"4a",x"bf",x"97",x"ff"),
   444 => (x"ea",x"c2",x"49",x"a1"),
   445 => (x"ea",x"c2",x"59",x"fe"),
   446 => (x"c5",x"49",x"bf",x"fa"),
   447 => (x"81",x"ff",x"c7",x"31"),
   448 => (x"ef",x"c2",x"29",x"c9"),
   449 => (x"e3",x"c2",x"59",x"d7"),
   450 => (x"4a",x"bf",x"97",x"c5"),
   451 => (x"e3",x"c2",x"32",x"c8"),
   452 => (x"4b",x"bf",x"97",x"c4"),
   453 => (x"66",x"c4",x"4a",x"a2"),
   454 => (x"c2",x"82",x"6e",x"92"),
   455 => (x"c2",x"5a",x"d3",x"ef"),
   456 => (x"c0",x"48",x"cb",x"ef"),
   457 => (x"c7",x"ef",x"c2",x"78"),
   458 => (x"78",x"a1",x"72",x"48"),
   459 => (x"48",x"d7",x"ef",x"c2"),
   460 => (x"bf",x"cb",x"ef",x"c2"),
   461 => (x"db",x"ef",x"c2",x"78"),
   462 => (x"cf",x"ef",x"c2",x"48"),
   463 => (x"ea",x"c2",x"78",x"bf"),
   464 => (x"c0",x"02",x"bf",x"f6"),
   465 => (x"48",x"74",x"87",x"c9"),
   466 => (x"7e",x"70",x"30",x"c4"),
   467 => (x"c2",x"87",x"c9",x"c0"),
   468 => (x"48",x"bf",x"d3",x"ef"),
   469 => (x"7e",x"70",x"30",x"c4"),
   470 => (x"48",x"fa",x"ea",x"c2"),
   471 => (x"48",x"c1",x"78",x"6e"),
   472 => (x"4d",x"26",x"8e",x"f8"),
   473 => (x"4b",x"26",x"4c",x"26"),
   474 => (x"5e",x"0e",x"4f",x"26"),
   475 => (x"0e",x"5d",x"5c",x"5b"),
   476 => (x"ea",x"c2",x"4a",x"71"),
   477 => (x"cb",x"02",x"bf",x"f6"),
   478 => (x"c7",x"4b",x"72",x"87"),
   479 => (x"c1",x"4c",x"72",x"2b"),
   480 => (x"87",x"c9",x"9c",x"ff"),
   481 => (x"2b",x"c8",x"4b",x"72"),
   482 => (x"ff",x"c3",x"4c",x"72"),
   483 => (x"c3",x"ef",x"c2",x"9c"),
   484 => (x"ef",x"c0",x"83",x"bf"),
   485 => (x"02",x"ab",x"bf",x"d0"),
   486 => (x"ef",x"c0",x"87",x"d9"),
   487 => (x"e2",x"c2",x"5b",x"d4"),
   488 => (x"49",x"73",x"1e",x"ee"),
   489 => (x"c4",x"87",x"fd",x"f0"),
   490 => (x"05",x"98",x"70",x"86"),
   491 => (x"48",x"c0",x"87",x"c5"),
   492 => (x"c2",x"87",x"e6",x"c0"),
   493 => (x"02",x"bf",x"f6",x"ea"),
   494 => (x"49",x"74",x"87",x"d2"),
   495 => (x"e2",x"c2",x"91",x"c4"),
   496 => (x"4d",x"69",x"81",x"ee"),
   497 => (x"ff",x"ff",x"ff",x"cf"),
   498 => (x"87",x"cb",x"9d",x"ff"),
   499 => (x"91",x"c2",x"49",x"74"),
   500 => (x"81",x"ee",x"e2",x"c2"),
   501 => (x"75",x"4d",x"69",x"9f"),
   502 => (x"87",x"c6",x"fe",x"48"),
   503 => (x"5c",x"5b",x"5e",x"0e"),
   504 => (x"86",x"f8",x"0e",x"5d"),
   505 => (x"05",x"9c",x"4c",x"71"),
   506 => (x"48",x"c0",x"87",x"c5"),
   507 => (x"c8",x"87",x"c2",x"c3"),
   508 => (x"48",x"6e",x"7e",x"a4"),
   509 => (x"66",x"d8",x"78",x"c0"),
   510 => (x"d8",x"87",x"c7",x"02"),
   511 => (x"05",x"bf",x"97",x"66"),
   512 => (x"48",x"c0",x"87",x"c5"),
   513 => (x"c0",x"87",x"ea",x"c2"),
   514 => (x"49",x"49",x"c1",x"1e"),
   515 => (x"c4",x"87",x"e6",x"c7"),
   516 => (x"9d",x"4d",x"70",x"86"),
   517 => (x"87",x"c2",x"c1",x"02"),
   518 => (x"4a",x"fe",x"ea",x"c2"),
   519 => (x"e0",x"49",x"66",x"d8"),
   520 => (x"98",x"70",x"87",x"ec"),
   521 => (x"87",x"f2",x"c0",x"02"),
   522 => (x"66",x"d8",x"4a",x"75"),
   523 => (x"e1",x"4b",x"cb",x"49"),
   524 => (x"98",x"70",x"87",x"d1"),
   525 => (x"87",x"e2",x"c0",x"02"),
   526 => (x"9d",x"75",x"1e",x"c0"),
   527 => (x"c8",x"87",x"c7",x"02"),
   528 => (x"78",x"c0",x"48",x"a6"),
   529 => (x"a6",x"c8",x"87",x"c5"),
   530 => (x"c8",x"78",x"c1",x"48"),
   531 => (x"e4",x"c6",x"49",x"66"),
   532 => (x"70",x"86",x"c4",x"87"),
   533 => (x"fe",x"05",x"9d",x"4d"),
   534 => (x"9d",x"75",x"87",x"fe"),
   535 => (x"87",x"cf",x"c1",x"02"),
   536 => (x"6e",x"49",x"a5",x"dc"),
   537 => (x"da",x"78",x"69",x"48"),
   538 => (x"a6",x"c4",x"49",x"a5"),
   539 => (x"78",x"a4",x"c4",x"48"),
   540 => (x"c4",x"48",x"69",x"9f"),
   541 => (x"c2",x"78",x"08",x"66"),
   542 => (x"02",x"bf",x"f6",x"ea"),
   543 => (x"a5",x"d4",x"87",x"d2"),
   544 => (x"49",x"69",x"9f",x"49"),
   545 => (x"99",x"ff",x"ff",x"c0"),
   546 => (x"30",x"d0",x"48",x"71"),
   547 => (x"87",x"c2",x"7e",x"70"),
   548 => (x"49",x"6e",x"7e",x"c0"),
   549 => (x"bf",x"66",x"c4",x"48"),
   550 => (x"08",x"66",x"c4",x"80"),
   551 => (x"cc",x"7c",x"c0",x"78"),
   552 => (x"66",x"c4",x"49",x"a4"),
   553 => (x"a4",x"d0",x"79",x"bf"),
   554 => (x"c1",x"79",x"c0",x"49"),
   555 => (x"c0",x"87",x"c2",x"48"),
   556 => (x"fa",x"8e",x"f8",x"48"),
   557 => (x"5e",x"0e",x"87",x"ec"),
   558 => (x"0e",x"5d",x"5c",x"5b"),
   559 => (x"02",x"9c",x"4c",x"71"),
   560 => (x"c8",x"87",x"ca",x"c1"),
   561 => (x"02",x"69",x"49",x"a4"),
   562 => (x"d0",x"87",x"c2",x"c1"),
   563 => (x"49",x"6c",x"4a",x"66"),
   564 => (x"5a",x"a6",x"d4",x"82"),
   565 => (x"b9",x"4d",x"66",x"d0"),
   566 => (x"bf",x"f2",x"ea",x"c2"),
   567 => (x"72",x"ba",x"ff",x"4a"),
   568 => (x"02",x"99",x"71",x"99"),
   569 => (x"c4",x"87",x"e4",x"c0"),
   570 => (x"49",x"6b",x"4b",x"a4"),
   571 => (x"70",x"87",x"fb",x"f9"),
   572 => (x"ee",x"ea",x"c2",x"7b"),
   573 => (x"81",x"6c",x"49",x"bf"),
   574 => (x"b9",x"75",x"7c",x"71"),
   575 => (x"bf",x"f2",x"ea",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"05",x"99",x"71",x"99"),
   578 => (x"75",x"87",x"dc",x"ff"),
   579 => (x"87",x"d2",x"f9",x"7c"),
   580 => (x"71",x"1e",x"73",x"1e"),
   581 => (x"c7",x"02",x"9b",x"4b"),
   582 => (x"49",x"a3",x"c8",x"87"),
   583 => (x"87",x"c5",x"05",x"69"),
   584 => (x"f7",x"c0",x"48",x"c0"),
   585 => (x"c7",x"ef",x"c2",x"87"),
   586 => (x"a3",x"c4",x"4a",x"bf"),
   587 => (x"c2",x"49",x"69",x"49"),
   588 => (x"ee",x"ea",x"c2",x"89"),
   589 => (x"a2",x"71",x"91",x"bf"),
   590 => (x"f2",x"ea",x"c2",x"4a"),
   591 => (x"99",x"6b",x"49",x"bf"),
   592 => (x"c0",x"4a",x"a2",x"71"),
   593 => (x"c8",x"5a",x"d4",x"ef"),
   594 => (x"49",x"72",x"1e",x"66"),
   595 => (x"c4",x"87",x"d5",x"ea"),
   596 => (x"05",x"98",x"70",x"86"),
   597 => (x"48",x"c0",x"87",x"c4"),
   598 => (x"48",x"c1",x"87",x"c2"),
   599 => (x"1e",x"87",x"c7",x"f8"),
   600 => (x"4b",x"71",x"1e",x"73"),
   601 => (x"e4",x"c0",x"02",x"9b"),
   602 => (x"db",x"ef",x"c2",x"87"),
   603 => (x"c2",x"4a",x"73",x"5b"),
   604 => (x"ee",x"ea",x"c2",x"8a"),
   605 => (x"c2",x"92",x"49",x"bf"),
   606 => (x"48",x"bf",x"c7",x"ef"),
   607 => (x"ef",x"c2",x"80",x"72"),
   608 => (x"48",x"71",x"58",x"df"),
   609 => (x"ea",x"c2",x"30",x"c4"),
   610 => (x"ed",x"c0",x"58",x"fe"),
   611 => (x"d7",x"ef",x"c2",x"87"),
   612 => (x"cb",x"ef",x"c2",x"48"),
   613 => (x"ef",x"c2",x"78",x"bf"),
   614 => (x"ef",x"c2",x"48",x"db"),
   615 => (x"c2",x"78",x"bf",x"cf"),
   616 => (x"02",x"bf",x"f6",x"ea"),
   617 => (x"ea",x"c2",x"87",x"c9"),
   618 => (x"c4",x"49",x"bf",x"ee"),
   619 => (x"c2",x"87",x"c7",x"31"),
   620 => (x"49",x"bf",x"d3",x"ef"),
   621 => (x"ea",x"c2",x"31",x"c4"),
   622 => (x"e9",x"f6",x"59",x"fe"),
   623 => (x"5b",x"5e",x"0e",x"87"),
   624 => (x"4a",x"71",x"0e",x"5c"),
   625 => (x"9a",x"72",x"4b",x"c0"),
   626 => (x"87",x"e1",x"c0",x"02"),
   627 => (x"9f",x"49",x"a2",x"da"),
   628 => (x"ea",x"c2",x"4b",x"69"),
   629 => (x"cf",x"02",x"bf",x"f6"),
   630 => (x"49",x"a2",x"d4",x"87"),
   631 => (x"4c",x"49",x"69",x"9f"),
   632 => (x"9c",x"ff",x"ff",x"c0"),
   633 => (x"87",x"c2",x"34",x"d0"),
   634 => (x"49",x"74",x"4c",x"c0"),
   635 => (x"fd",x"49",x"73",x"b3"),
   636 => (x"ef",x"f5",x"87",x"ed"),
   637 => (x"5b",x"5e",x"0e",x"87"),
   638 => (x"f4",x"0e",x"5d",x"5c"),
   639 => (x"c0",x"4a",x"71",x"86"),
   640 => (x"02",x"9a",x"72",x"7e"),
   641 => (x"e2",x"c2",x"87",x"d8"),
   642 => (x"78",x"c0",x"48",x"ea"),
   643 => (x"48",x"e2",x"e2",x"c2"),
   644 => (x"bf",x"db",x"ef",x"c2"),
   645 => (x"e6",x"e2",x"c2",x"78"),
   646 => (x"d7",x"ef",x"c2",x"48"),
   647 => (x"eb",x"c2",x"78",x"bf"),
   648 => (x"50",x"c0",x"48",x"cb"),
   649 => (x"bf",x"fa",x"ea",x"c2"),
   650 => (x"ea",x"e2",x"c2",x"49"),
   651 => (x"aa",x"71",x"4a",x"bf"),
   652 => (x"87",x"c9",x"c4",x"03"),
   653 => (x"99",x"cf",x"49",x"72"),
   654 => (x"87",x"e9",x"c0",x"05"),
   655 => (x"48",x"d0",x"ef",x"c0"),
   656 => (x"bf",x"e2",x"e2",x"c2"),
   657 => (x"ee",x"e2",x"c2",x"78"),
   658 => (x"e2",x"e2",x"c2",x"1e"),
   659 => (x"e2",x"c2",x"49",x"bf"),
   660 => (x"a1",x"c1",x"48",x"e2"),
   661 => (x"cb",x"e6",x"71",x"78"),
   662 => (x"c0",x"86",x"c4",x"87"),
   663 => (x"c2",x"48",x"cc",x"ef"),
   664 => (x"cc",x"78",x"ee",x"e2"),
   665 => (x"cc",x"ef",x"c0",x"87"),
   666 => (x"e0",x"c0",x"48",x"bf"),
   667 => (x"d0",x"ef",x"c0",x"80"),
   668 => (x"ea",x"e2",x"c2",x"58"),
   669 => (x"80",x"c1",x"48",x"bf"),
   670 => (x"58",x"ee",x"e2",x"c2"),
   671 => (x"00",x"0b",x"cc",x"27"),
   672 => (x"bf",x"97",x"bf",x"00"),
   673 => (x"c2",x"02",x"9d",x"4d"),
   674 => (x"e5",x"c3",x"87",x"e3"),
   675 => (x"dc",x"c2",x"02",x"ad"),
   676 => (x"cc",x"ef",x"c0",x"87"),
   677 => (x"a3",x"cb",x"4b",x"bf"),
   678 => (x"cf",x"4c",x"11",x"49"),
   679 => (x"d2",x"c1",x"05",x"ac"),
   680 => (x"df",x"49",x"75",x"87"),
   681 => (x"cd",x"89",x"c1",x"99"),
   682 => (x"fe",x"ea",x"c2",x"91"),
   683 => (x"4a",x"a3",x"c1",x"81"),
   684 => (x"a3",x"c3",x"51",x"12"),
   685 => (x"c5",x"51",x"12",x"4a"),
   686 => (x"51",x"12",x"4a",x"a3"),
   687 => (x"12",x"4a",x"a3",x"c7"),
   688 => (x"4a",x"a3",x"c9",x"51"),
   689 => (x"a3",x"ce",x"51",x"12"),
   690 => (x"d0",x"51",x"12",x"4a"),
   691 => (x"51",x"12",x"4a",x"a3"),
   692 => (x"12",x"4a",x"a3",x"d2"),
   693 => (x"4a",x"a3",x"d4",x"51"),
   694 => (x"a3",x"d6",x"51",x"12"),
   695 => (x"d8",x"51",x"12",x"4a"),
   696 => (x"51",x"12",x"4a",x"a3"),
   697 => (x"12",x"4a",x"a3",x"dc"),
   698 => (x"4a",x"a3",x"de",x"51"),
   699 => (x"7e",x"c1",x"51",x"12"),
   700 => (x"74",x"87",x"fa",x"c0"),
   701 => (x"05",x"99",x"c8",x"49"),
   702 => (x"74",x"87",x"eb",x"c0"),
   703 => (x"05",x"99",x"d0",x"49"),
   704 => (x"66",x"dc",x"87",x"d1"),
   705 => (x"87",x"cb",x"c0",x"02"),
   706 => (x"66",x"dc",x"49",x"73"),
   707 => (x"02",x"98",x"70",x"0f"),
   708 => (x"6e",x"87",x"d3",x"c0"),
   709 => (x"87",x"c6",x"c0",x"05"),
   710 => (x"48",x"fe",x"ea",x"c2"),
   711 => (x"ef",x"c0",x"50",x"c0"),
   712 => (x"c2",x"48",x"bf",x"cc"),
   713 => (x"eb",x"c2",x"87",x"e1"),
   714 => (x"50",x"c0",x"48",x"cb"),
   715 => (x"fa",x"ea",x"c2",x"7e"),
   716 => (x"e2",x"c2",x"49",x"bf"),
   717 => (x"71",x"4a",x"bf",x"ea"),
   718 => (x"f7",x"fb",x"04",x"aa"),
   719 => (x"db",x"ef",x"c2",x"87"),
   720 => (x"c8",x"c0",x"05",x"bf"),
   721 => (x"f6",x"ea",x"c2",x"87"),
   722 => (x"f8",x"c1",x"02",x"bf"),
   723 => (x"e6",x"e2",x"c2",x"87"),
   724 => (x"d5",x"f0",x"49",x"bf"),
   725 => (x"c2",x"49",x"70",x"87"),
   726 => (x"c4",x"59",x"ea",x"e2"),
   727 => (x"e2",x"c2",x"48",x"a6"),
   728 => (x"c2",x"78",x"bf",x"e6"),
   729 => (x"02",x"bf",x"f6",x"ea"),
   730 => (x"c4",x"87",x"d8",x"c0"),
   731 => (x"ff",x"cf",x"49",x"66"),
   732 => (x"99",x"f8",x"ff",x"ff"),
   733 => (x"c5",x"c0",x"02",x"a9"),
   734 => (x"c0",x"4c",x"c0",x"87"),
   735 => (x"4c",x"c1",x"87",x"e1"),
   736 => (x"c4",x"87",x"dc",x"c0"),
   737 => (x"ff",x"cf",x"49",x"66"),
   738 => (x"02",x"a9",x"99",x"f8"),
   739 => (x"c8",x"87",x"c8",x"c0"),
   740 => (x"78",x"c0",x"48",x"a6"),
   741 => (x"c8",x"87",x"c5",x"c0"),
   742 => (x"78",x"c1",x"48",x"a6"),
   743 => (x"74",x"4c",x"66",x"c8"),
   744 => (x"e0",x"c0",x"05",x"9c"),
   745 => (x"49",x"66",x"c4",x"87"),
   746 => (x"ea",x"c2",x"89",x"c2"),
   747 => (x"91",x"4a",x"bf",x"ee"),
   748 => (x"bf",x"c7",x"ef",x"c2"),
   749 => (x"e2",x"e2",x"c2",x"4a"),
   750 => (x"78",x"a1",x"72",x"48"),
   751 => (x"48",x"ea",x"e2",x"c2"),
   752 => (x"df",x"f9",x"78",x"c0"),
   753 => (x"f4",x"48",x"c0",x"87"),
   754 => (x"87",x"d6",x"ee",x"8e"),
   755 => (x"00",x"00",x"00",x"00"),
   756 => (x"ff",x"ff",x"ff",x"ff"),
   757 => (x"00",x"00",x"0b",x"dc"),
   758 => (x"00",x"00",x"0b",x"e5"),
   759 => (x"33",x"54",x"41",x"46"),
   760 => (x"20",x"20",x"20",x"32"),
   761 => (x"54",x"41",x"46",x"00"),
   762 => (x"20",x"20",x"36",x"31"),
   763 => (x"ff",x"1e",x"00",x"20"),
   764 => (x"ff",x"c3",x"48",x"d4"),
   765 => (x"26",x"48",x"68",x"78"),
   766 => (x"d4",x"ff",x"1e",x"4f"),
   767 => (x"78",x"ff",x"c3",x"48"),
   768 => (x"c0",x"48",x"d0",x"ff"),
   769 => (x"d4",x"ff",x"78",x"e1"),
   770 => (x"c2",x"78",x"d4",x"48"),
   771 => (x"ff",x"48",x"df",x"ef"),
   772 => (x"26",x"50",x"bf",x"d4"),
   773 => (x"d0",x"ff",x"1e",x"4f"),
   774 => (x"78",x"e0",x"c0",x"48"),
   775 => (x"ff",x"1e",x"4f",x"26"),
   776 => (x"49",x"70",x"87",x"cc"),
   777 => (x"87",x"c6",x"02",x"99"),
   778 => (x"05",x"a9",x"fb",x"c0"),
   779 => (x"48",x"71",x"87",x"f1"),
   780 => (x"5e",x"0e",x"4f",x"26"),
   781 => (x"71",x"0e",x"5c",x"5b"),
   782 => (x"fe",x"4c",x"c0",x"4b"),
   783 => (x"49",x"70",x"87",x"f0"),
   784 => (x"f9",x"c0",x"02",x"99"),
   785 => (x"a9",x"ec",x"c0",x"87"),
   786 => (x"87",x"f2",x"c0",x"02"),
   787 => (x"02",x"a9",x"fb",x"c0"),
   788 => (x"cc",x"87",x"eb",x"c0"),
   789 => (x"03",x"ac",x"b7",x"66"),
   790 => (x"66",x"d0",x"87",x"c7"),
   791 => (x"71",x"87",x"c2",x"02"),
   792 => (x"02",x"99",x"71",x"53"),
   793 => (x"84",x"c1",x"87",x"c2"),
   794 => (x"70",x"87",x"c3",x"fe"),
   795 => (x"cd",x"02",x"99",x"49"),
   796 => (x"a9",x"ec",x"c0",x"87"),
   797 => (x"c0",x"87",x"c7",x"02"),
   798 => (x"ff",x"05",x"a9",x"fb"),
   799 => (x"66",x"d0",x"87",x"d5"),
   800 => (x"c0",x"87",x"c3",x"02"),
   801 => (x"ec",x"c0",x"7b",x"97"),
   802 => (x"87",x"c4",x"05",x"a9"),
   803 => (x"87",x"c5",x"4a",x"74"),
   804 => (x"0a",x"c0",x"4a",x"74"),
   805 => (x"c2",x"48",x"72",x"8a"),
   806 => (x"26",x"4d",x"26",x"87"),
   807 => (x"26",x"4b",x"26",x"4c"),
   808 => (x"c9",x"fd",x"1e",x"4f"),
   809 => (x"4a",x"49",x"70",x"87"),
   810 => (x"04",x"aa",x"f0",x"c0"),
   811 => (x"f9",x"c0",x"87",x"c9"),
   812 => (x"87",x"c3",x"01",x"aa"),
   813 => (x"c1",x"8a",x"f0",x"c0"),
   814 => (x"c9",x"04",x"aa",x"c1"),
   815 => (x"aa",x"da",x"c1",x"87"),
   816 => (x"c0",x"87",x"c3",x"01"),
   817 => (x"48",x"72",x"8a",x"f7"),
   818 => (x"5e",x"0e",x"4f",x"26"),
   819 => (x"71",x"0e",x"5c",x"5b"),
   820 => (x"4b",x"d4",x"ff",x"4a"),
   821 => (x"e7",x"c0",x"49",x"72"),
   822 => (x"9c",x"4c",x"70",x"87"),
   823 => (x"c1",x"87",x"c2",x"02"),
   824 => (x"48",x"d0",x"ff",x"8c"),
   825 => (x"d5",x"c1",x"78",x"c5"),
   826 => (x"c6",x"49",x"74",x"7b"),
   827 => (x"fc",x"e0",x"c1",x"31"),
   828 => (x"48",x"4a",x"bf",x"97"),
   829 => (x"7b",x"70",x"b0",x"71"),
   830 => (x"c4",x"48",x"d0",x"ff"),
   831 => (x"87",x"db",x"fe",x"78"),
   832 => (x"5c",x"5b",x"5e",x"0e"),
   833 => (x"86",x"f8",x"0e",x"5d"),
   834 => (x"7e",x"c0",x"4c",x"71"),
   835 => (x"c0",x"87",x"ea",x"fb"),
   836 => (x"ed",x"f6",x"c0",x"4b"),
   837 => (x"c0",x"49",x"bf",x"97"),
   838 => (x"87",x"cf",x"04",x"a9"),
   839 => (x"c1",x"87",x"ff",x"fb"),
   840 => (x"ed",x"f6",x"c0",x"83"),
   841 => (x"ab",x"49",x"bf",x"97"),
   842 => (x"c0",x"87",x"f1",x"06"),
   843 => (x"bf",x"97",x"ed",x"f6"),
   844 => (x"fa",x"87",x"cf",x"02"),
   845 => (x"49",x"70",x"87",x"f8"),
   846 => (x"87",x"c6",x"02",x"99"),
   847 => (x"05",x"a9",x"ec",x"c0"),
   848 => (x"4b",x"c0",x"87",x"f1"),
   849 => (x"70",x"87",x"e7",x"fa"),
   850 => (x"87",x"e2",x"fa",x"4d"),
   851 => (x"fa",x"58",x"a6",x"c8"),
   852 => (x"4a",x"70",x"87",x"dc"),
   853 => (x"a4",x"c8",x"83",x"c1"),
   854 => (x"49",x"69",x"97",x"49"),
   855 => (x"87",x"c7",x"02",x"ad"),
   856 => (x"05",x"ad",x"ff",x"c0"),
   857 => (x"c9",x"87",x"e7",x"c0"),
   858 => (x"69",x"97",x"49",x"a4"),
   859 => (x"a9",x"66",x"c4",x"49"),
   860 => (x"48",x"87",x"c7",x"02"),
   861 => (x"05",x"a8",x"ff",x"c0"),
   862 => (x"a4",x"ca",x"87",x"d4"),
   863 => (x"49",x"69",x"97",x"49"),
   864 => (x"87",x"c6",x"02",x"aa"),
   865 => (x"05",x"aa",x"ff",x"c0"),
   866 => (x"7e",x"c1",x"87",x"c4"),
   867 => (x"ec",x"c0",x"87",x"d0"),
   868 => (x"87",x"c6",x"02",x"ad"),
   869 => (x"05",x"ad",x"fb",x"c0"),
   870 => (x"4b",x"c0",x"87",x"c4"),
   871 => (x"02",x"6e",x"7e",x"c1"),
   872 => (x"f9",x"87",x"e1",x"fe"),
   873 => (x"48",x"73",x"87",x"ef"),
   874 => (x"ec",x"fb",x"8e",x"f8"),
   875 => (x"5e",x"0e",x"00",x"87"),
   876 => (x"0e",x"5d",x"5c",x"5b"),
   877 => (x"4d",x"71",x"86",x"f8"),
   878 => (x"75",x"4b",x"d4",x"ff"),
   879 => (x"e4",x"ef",x"c2",x"1e"),
   880 => (x"87",x"d8",x"e8",x"49"),
   881 => (x"98",x"70",x"86",x"c4"),
   882 => (x"87",x"cc",x"c4",x"02"),
   883 => (x"c1",x"48",x"a6",x"c4"),
   884 => (x"78",x"bf",x"fe",x"e0"),
   885 => (x"f1",x"fb",x"49",x"75"),
   886 => (x"48",x"d0",x"ff",x"87"),
   887 => (x"d6",x"c1",x"78",x"c5"),
   888 => (x"75",x"4a",x"c0",x"7b"),
   889 => (x"7b",x"11",x"49",x"a2"),
   890 => (x"b7",x"cb",x"82",x"c1"),
   891 => (x"87",x"f3",x"04",x"aa"),
   892 => (x"ff",x"c3",x"4a",x"cc"),
   893 => (x"c0",x"82",x"c1",x"7b"),
   894 => (x"04",x"aa",x"b7",x"e0"),
   895 => (x"d0",x"ff",x"87",x"f4"),
   896 => (x"c3",x"78",x"c4",x"48"),
   897 => (x"78",x"c5",x"7b",x"ff"),
   898 => (x"c1",x"7b",x"d3",x"c1"),
   899 => (x"66",x"78",x"c4",x"7b"),
   900 => (x"a8",x"b7",x"c0",x"48"),
   901 => (x"87",x"f0",x"c2",x"06"),
   902 => (x"bf",x"ec",x"ef",x"c2"),
   903 => (x"48",x"66",x"c4",x"4c"),
   904 => (x"a6",x"c8",x"88",x"74"),
   905 => (x"02",x"9c",x"74",x"58"),
   906 => (x"c2",x"87",x"f9",x"c1"),
   907 => (x"c8",x"7e",x"ee",x"e2"),
   908 => (x"c0",x"8c",x"4d",x"c0"),
   909 => (x"c6",x"03",x"ac",x"b7"),
   910 => (x"a4",x"c0",x"c8",x"87"),
   911 => (x"c2",x"4c",x"c0",x"4d"),
   912 => (x"bf",x"97",x"df",x"ef"),
   913 => (x"02",x"99",x"d0",x"49"),
   914 => (x"1e",x"c0",x"87",x"d1"),
   915 => (x"49",x"e4",x"ef",x"c2"),
   916 => (x"c4",x"87",x"fd",x"ea"),
   917 => (x"4a",x"49",x"70",x"86"),
   918 => (x"c2",x"87",x"ee",x"c0"),
   919 => (x"c2",x"1e",x"ee",x"e2"),
   920 => (x"ea",x"49",x"e4",x"ef"),
   921 => (x"86",x"c4",x"87",x"ea"),
   922 => (x"ff",x"4a",x"49",x"70"),
   923 => (x"c5",x"c8",x"48",x"d0"),
   924 => (x"7b",x"d4",x"c1",x"78"),
   925 => (x"7b",x"bf",x"97",x"6e"),
   926 => (x"80",x"c1",x"48",x"6e"),
   927 => (x"8d",x"c1",x"7e",x"70"),
   928 => (x"87",x"f0",x"ff",x"05"),
   929 => (x"c4",x"48",x"d0",x"ff"),
   930 => (x"05",x"9a",x"72",x"78"),
   931 => (x"48",x"c0",x"87",x"c5"),
   932 => (x"c1",x"87",x"c7",x"c1"),
   933 => (x"e4",x"ef",x"c2",x"1e"),
   934 => (x"87",x"da",x"e8",x"49"),
   935 => (x"9c",x"74",x"86",x"c4"),
   936 => (x"87",x"c7",x"fe",x"05"),
   937 => (x"c0",x"48",x"66",x"c4"),
   938 => (x"d1",x"06",x"a8",x"b7"),
   939 => (x"e4",x"ef",x"c2",x"87"),
   940 => (x"d0",x"78",x"c0",x"48"),
   941 => (x"f4",x"78",x"c0",x"80"),
   942 => (x"f0",x"ef",x"c2",x"80"),
   943 => (x"66",x"c4",x"78",x"bf"),
   944 => (x"a8",x"b7",x"c0",x"48"),
   945 => (x"87",x"d0",x"fd",x"01"),
   946 => (x"c5",x"48",x"d0",x"ff"),
   947 => (x"7b",x"d3",x"c1",x"78"),
   948 => (x"78",x"c4",x"7b",x"c0"),
   949 => (x"87",x"c2",x"48",x"c1"),
   950 => (x"8e",x"f8",x"48",x"c0"),
   951 => (x"4c",x"26",x"4d",x"26"),
   952 => (x"4f",x"26",x"4b",x"26"),
   953 => (x"5c",x"5b",x"5e",x"0e"),
   954 => (x"71",x"1e",x"0e",x"5d"),
   955 => (x"4d",x"4c",x"c0",x"4b"),
   956 => (x"e8",x"c0",x"04",x"ab"),
   957 => (x"c0",x"f4",x"c0",x"87"),
   958 => (x"02",x"9d",x"75",x"1e"),
   959 => (x"4a",x"c0",x"87",x"c4"),
   960 => (x"4a",x"c1",x"87",x"c2"),
   961 => (x"ec",x"eb",x"49",x"72"),
   962 => (x"70",x"86",x"c4",x"87"),
   963 => (x"6e",x"84",x"c1",x"7e"),
   964 => (x"73",x"87",x"c2",x"05"),
   965 => (x"73",x"85",x"c1",x"4c"),
   966 => (x"d8",x"ff",x"06",x"ac"),
   967 => (x"26",x"48",x"6e",x"87"),
   968 => (x"1e",x"87",x"f9",x"fe"),
   969 => (x"66",x"c4",x"4a",x"71"),
   970 => (x"72",x"87",x"c5",x"05"),
   971 => (x"87",x"fe",x"f9",x"49"),
   972 => (x"5e",x"0e",x"4f",x"26"),
   973 => (x"0e",x"5d",x"5c",x"5b"),
   974 => (x"49",x"4c",x"71",x"1e"),
   975 => (x"f0",x"c2",x"91",x"de"),
   976 => (x"85",x"71",x"4d",x"cc"),
   977 => (x"c1",x"02",x"6d",x"97"),
   978 => (x"ef",x"c2",x"87",x"dd"),
   979 => (x"74",x"4a",x"bf",x"f8"),
   980 => (x"fe",x"49",x"72",x"82"),
   981 => (x"7e",x"70",x"87",x"ce"),
   982 => (x"c0",x"02",x"98",x"48"),
   983 => (x"f0",x"c2",x"87",x"f2"),
   984 => (x"4a",x"70",x"4b",x"c0"),
   985 => (x"c4",x"ff",x"49",x"cb"),
   986 => (x"4b",x"74",x"87",x"fd"),
   987 => (x"e1",x"c1",x"93",x"cb"),
   988 => (x"83",x"c4",x"83",x"d0"),
   989 => (x"7b",x"eb",x"fe",x"c0"),
   990 => (x"c1",x"c1",x"49",x"74"),
   991 => (x"7b",x"75",x"87",x"f3"),
   992 => (x"97",x"fd",x"e0",x"c1"),
   993 => (x"c2",x"1e",x"49",x"bf"),
   994 => (x"fe",x"49",x"c0",x"f0"),
   995 => (x"86",x"c4",x"87",x"d5"),
   996 => (x"c1",x"c1",x"49",x"74"),
   997 => (x"49",x"c0",x"87",x"db"),
   998 => (x"87",x"fa",x"c2",x"c1"),
   999 => (x"48",x"e0",x"ef",x"c2"),
  1000 => (x"49",x"c1",x"78",x"c0"),
  1001 => (x"26",x"87",x"dc",x"de"),
  1002 => (x"4c",x"87",x"f1",x"fc"),
  1003 => (x"69",x"64",x"61",x"6f"),
  1004 => (x"2e",x"2e",x"67",x"6e"),
  1005 => (x"5e",x"0e",x"00",x"2e"),
  1006 => (x"71",x"0e",x"5c",x"5b"),
  1007 => (x"ef",x"c2",x"4a",x"4b"),
  1008 => (x"72",x"82",x"bf",x"f8"),
  1009 => (x"87",x"dc",x"fc",x"49"),
  1010 => (x"02",x"9c",x"4c",x"70"),
  1011 => (x"e7",x"49",x"87",x"c4"),
  1012 => (x"ef",x"c2",x"87",x"eb"),
  1013 => (x"78",x"c0",x"48",x"f8"),
  1014 => (x"e6",x"dd",x"49",x"c1"),
  1015 => (x"87",x"fe",x"fb",x"87"),
  1016 => (x"5c",x"5b",x"5e",x"0e"),
  1017 => (x"86",x"f4",x"0e",x"5d"),
  1018 => (x"4d",x"ee",x"e2",x"c2"),
  1019 => (x"a6",x"c4",x"4c",x"c0"),
  1020 => (x"c2",x"78",x"c0",x"48"),
  1021 => (x"49",x"bf",x"f8",x"ef"),
  1022 => (x"c1",x"06",x"a9",x"c0"),
  1023 => (x"e2",x"c2",x"87",x"c1"),
  1024 => (x"02",x"98",x"48",x"ee"),
  1025 => (x"c0",x"87",x"f8",x"c0"),
  1026 => (x"c8",x"1e",x"c0",x"f4"),
  1027 => (x"87",x"c7",x"02",x"66"),
  1028 => (x"c0",x"48",x"a6",x"c4"),
  1029 => (x"c4",x"87",x"c5",x"78"),
  1030 => (x"78",x"c1",x"48",x"a6"),
  1031 => (x"e7",x"49",x"66",x"c4"),
  1032 => (x"86",x"c4",x"87",x"d3"),
  1033 => (x"84",x"c1",x"4d",x"70"),
  1034 => (x"c1",x"48",x"66",x"c4"),
  1035 => (x"58",x"a6",x"c8",x"80"),
  1036 => (x"bf",x"f8",x"ef",x"c2"),
  1037 => (x"c6",x"03",x"ac",x"49"),
  1038 => (x"05",x"9d",x"75",x"87"),
  1039 => (x"c0",x"87",x"c8",x"ff"),
  1040 => (x"02",x"9d",x"75",x"4c"),
  1041 => (x"c0",x"87",x"e0",x"c3"),
  1042 => (x"c8",x"1e",x"c0",x"f4"),
  1043 => (x"87",x"c7",x"02",x"66"),
  1044 => (x"c0",x"48",x"a6",x"cc"),
  1045 => (x"cc",x"87",x"c5",x"78"),
  1046 => (x"78",x"c1",x"48",x"a6"),
  1047 => (x"e6",x"49",x"66",x"cc"),
  1048 => (x"86",x"c4",x"87",x"d3"),
  1049 => (x"98",x"48",x"7e",x"70"),
  1050 => (x"87",x"e8",x"c2",x"02"),
  1051 => (x"97",x"81",x"cb",x"49"),
  1052 => (x"99",x"d0",x"49",x"69"),
  1053 => (x"87",x"d6",x"c1",x"02"),
  1054 => (x"4a",x"f6",x"fe",x"c0"),
  1055 => (x"91",x"cb",x"49",x"74"),
  1056 => (x"81",x"d0",x"e1",x"c1"),
  1057 => (x"81",x"c8",x"79",x"72"),
  1058 => (x"74",x"51",x"ff",x"c3"),
  1059 => (x"c2",x"91",x"de",x"49"),
  1060 => (x"71",x"4d",x"cc",x"f0"),
  1061 => (x"97",x"c1",x"c2",x"85"),
  1062 => (x"49",x"a5",x"c1",x"7d"),
  1063 => (x"c2",x"51",x"e0",x"c0"),
  1064 => (x"bf",x"97",x"fe",x"ea"),
  1065 => (x"c1",x"87",x"d2",x"02"),
  1066 => (x"4b",x"a5",x"c2",x"84"),
  1067 => (x"4a",x"fe",x"ea",x"c2"),
  1068 => (x"ff",x"fe",x"49",x"db"),
  1069 => (x"db",x"c1",x"87",x"f1"),
  1070 => (x"49",x"a5",x"cd",x"87"),
  1071 => (x"84",x"c1",x"51",x"c0"),
  1072 => (x"6e",x"4b",x"a5",x"c2"),
  1073 => (x"fe",x"49",x"cb",x"4a"),
  1074 => (x"c1",x"87",x"dc",x"ff"),
  1075 => (x"fc",x"c0",x"87",x"c6"),
  1076 => (x"49",x"74",x"4a",x"f2"),
  1077 => (x"e1",x"c1",x"91",x"cb"),
  1078 => (x"79",x"72",x"81",x"d0"),
  1079 => (x"97",x"fe",x"ea",x"c2"),
  1080 => (x"87",x"d8",x"02",x"bf"),
  1081 => (x"91",x"de",x"49",x"74"),
  1082 => (x"f0",x"c2",x"84",x"c1"),
  1083 => (x"83",x"71",x"4b",x"cc"),
  1084 => (x"4a",x"fe",x"ea",x"c2"),
  1085 => (x"fe",x"fe",x"49",x"dd"),
  1086 => (x"87",x"d8",x"87",x"ed"),
  1087 => (x"93",x"de",x"4b",x"74"),
  1088 => (x"83",x"cc",x"f0",x"c2"),
  1089 => (x"c0",x"49",x"a3",x"cb"),
  1090 => (x"73",x"84",x"c1",x"51"),
  1091 => (x"49",x"cb",x"4a",x"6e"),
  1092 => (x"87",x"d3",x"fe",x"fe"),
  1093 => (x"c1",x"48",x"66",x"c4"),
  1094 => (x"58",x"a6",x"c8",x"80"),
  1095 => (x"c0",x"03",x"ac",x"c7"),
  1096 => (x"05",x"6e",x"87",x"c5"),
  1097 => (x"74",x"87",x"e0",x"fc"),
  1098 => (x"f6",x"8e",x"f4",x"48"),
  1099 => (x"73",x"1e",x"87",x"ee"),
  1100 => (x"49",x"4b",x"71",x"1e"),
  1101 => (x"e1",x"c1",x"91",x"cb"),
  1102 => (x"a1",x"c8",x"81",x"d0"),
  1103 => (x"fc",x"e0",x"c1",x"4a"),
  1104 => (x"c9",x"50",x"12",x"48"),
  1105 => (x"f6",x"c0",x"4a",x"a1"),
  1106 => (x"50",x"12",x"48",x"ed"),
  1107 => (x"e0",x"c1",x"81",x"ca"),
  1108 => (x"50",x"11",x"48",x"fd"),
  1109 => (x"97",x"fd",x"e0",x"c1"),
  1110 => (x"c0",x"1e",x"49",x"bf"),
  1111 => (x"87",x"c3",x"f7",x"49"),
  1112 => (x"48",x"e0",x"ef",x"c2"),
  1113 => (x"49",x"c1",x"78",x"de"),
  1114 => (x"26",x"87",x"d8",x"d7"),
  1115 => (x"1e",x"87",x"f1",x"f5"),
  1116 => (x"cb",x"49",x"4a",x"71"),
  1117 => (x"d0",x"e1",x"c1",x"91"),
  1118 => (x"11",x"81",x"c8",x"81"),
  1119 => (x"e4",x"ef",x"c2",x"48"),
  1120 => (x"f8",x"ef",x"c2",x"58"),
  1121 => (x"c1",x"78",x"c0",x"48"),
  1122 => (x"87",x"f7",x"d6",x"49"),
  1123 => (x"c0",x"1e",x"4f",x"26"),
  1124 => (x"c1",x"fb",x"c0",x"49"),
  1125 => (x"1e",x"4f",x"26",x"87"),
  1126 => (x"d2",x"02",x"99",x"71"),
  1127 => (x"e5",x"e2",x"c1",x"87"),
  1128 => (x"f7",x"50",x"c0",x"48"),
  1129 => (x"ef",x"c5",x"c1",x"80"),
  1130 => (x"c9",x"e1",x"c1",x"40"),
  1131 => (x"c1",x"87",x"ce",x"78"),
  1132 => (x"c1",x"48",x"e1",x"e2"),
  1133 => (x"fc",x"78",x"c2",x"e1"),
  1134 => (x"ce",x"c6",x"c1",x"80"),
  1135 => (x"0e",x"4f",x"26",x"78"),
  1136 => (x"5d",x"5c",x"5b",x"5e"),
  1137 => (x"71",x"86",x"f4",x"0e"),
  1138 => (x"91",x"cb",x"49",x"4d"),
  1139 => (x"81",x"d0",x"e1",x"c1"),
  1140 => (x"ca",x"4a",x"a1",x"c8"),
  1141 => (x"a6",x"c4",x"7e",x"a1"),
  1142 => (x"e8",x"f3",x"c2",x"48"),
  1143 => (x"97",x"6e",x"78",x"bf"),
  1144 => (x"66",x"c4",x"4b",x"bf"),
  1145 => (x"70",x"28",x"73",x"48"),
  1146 => (x"48",x"12",x"4c",x"4b"),
  1147 => (x"70",x"58",x"a6",x"cc"),
  1148 => (x"c9",x"84",x"c1",x"9c"),
  1149 => (x"49",x"69",x"97",x"81"),
  1150 => (x"c2",x"04",x"ac",x"b7"),
  1151 => (x"6e",x"4c",x"c0",x"87"),
  1152 => (x"c8",x"4a",x"bf",x"97"),
  1153 => (x"31",x"72",x"49",x"66"),
  1154 => (x"66",x"c4",x"b9",x"ff"),
  1155 => (x"72",x"48",x"74",x"99"),
  1156 => (x"48",x"4a",x"70",x"30"),
  1157 => (x"f3",x"c2",x"b0",x"71"),
  1158 => (x"e5",x"c0",x"58",x"ec"),
  1159 => (x"49",x"c0",x"87",x"d3"),
  1160 => (x"75",x"87",x"e0",x"d4"),
  1161 => (x"c8",x"f7",x"c0",x"49"),
  1162 => (x"f2",x"8e",x"f4",x"87"),
  1163 => (x"73",x"1e",x"87",x"ee"),
  1164 => (x"49",x"4b",x"71",x"1e"),
  1165 => (x"73",x"87",x"c8",x"fe"),
  1166 => (x"87",x"c3",x"fe",x"49"),
  1167 => (x"1e",x"87",x"e1",x"f2"),
  1168 => (x"4b",x"71",x"1e",x"73"),
  1169 => (x"02",x"4a",x"a3",x"c6"),
  1170 => (x"8a",x"c1",x"87",x"db"),
  1171 => (x"8a",x"87",x"d6",x"02"),
  1172 => (x"87",x"da",x"c1",x"02"),
  1173 => (x"fc",x"c0",x"02",x"8a"),
  1174 => (x"c0",x"02",x"8a",x"87"),
  1175 => (x"02",x"8a",x"87",x"e1"),
  1176 => (x"db",x"c1",x"87",x"cb"),
  1177 => (x"fc",x"49",x"c7",x"87"),
  1178 => (x"de",x"c1",x"87",x"c5"),
  1179 => (x"f8",x"ef",x"c2",x"87"),
  1180 => (x"cb",x"c1",x"02",x"bf"),
  1181 => (x"88",x"c1",x"48",x"87"),
  1182 => (x"58",x"fc",x"ef",x"c2"),
  1183 => (x"c2",x"87",x"c1",x"c1"),
  1184 => (x"02",x"bf",x"fc",x"ef"),
  1185 => (x"c2",x"87",x"f9",x"c0"),
  1186 => (x"48",x"bf",x"f8",x"ef"),
  1187 => (x"ef",x"c2",x"80",x"c1"),
  1188 => (x"eb",x"c0",x"58",x"fc"),
  1189 => (x"f8",x"ef",x"c2",x"87"),
  1190 => (x"89",x"c6",x"49",x"bf"),
  1191 => (x"59",x"fc",x"ef",x"c2"),
  1192 => (x"03",x"a9",x"b7",x"c0"),
  1193 => (x"ef",x"c2",x"87",x"da"),
  1194 => (x"78",x"c0",x"48",x"f8"),
  1195 => (x"ef",x"c2",x"87",x"d2"),
  1196 => (x"cb",x"02",x"bf",x"fc"),
  1197 => (x"f8",x"ef",x"c2",x"87"),
  1198 => (x"80",x"c6",x"48",x"bf"),
  1199 => (x"58",x"fc",x"ef",x"c2"),
  1200 => (x"fe",x"d1",x"49",x"c0"),
  1201 => (x"c0",x"49",x"73",x"87"),
  1202 => (x"f0",x"87",x"e6",x"f4"),
  1203 => (x"5e",x"0e",x"87",x"d2"),
  1204 => (x"0e",x"5d",x"5c",x"5b"),
  1205 => (x"dc",x"86",x"d0",x"ff"),
  1206 => (x"a6",x"c8",x"59",x"a6"),
  1207 => (x"c4",x"78",x"c0",x"48"),
  1208 => (x"66",x"c4",x"c1",x"80"),
  1209 => (x"c1",x"80",x"c4",x"78"),
  1210 => (x"c1",x"80",x"c4",x"78"),
  1211 => (x"fc",x"ef",x"c2",x"78"),
  1212 => (x"c2",x"78",x"c1",x"48"),
  1213 => (x"48",x"bf",x"e0",x"ef"),
  1214 => (x"cb",x"05",x"a8",x"de"),
  1215 => (x"87",x"e0",x"f3",x"87"),
  1216 => (x"a6",x"cc",x"49",x"70"),
  1217 => (x"87",x"fa",x"cf",x"59"),
  1218 => (x"e4",x"87",x"ee",x"e3"),
  1219 => (x"dd",x"e3",x"87",x"d0"),
  1220 => (x"c0",x"4c",x"70",x"87"),
  1221 => (x"c1",x"02",x"ac",x"fb"),
  1222 => (x"66",x"d8",x"87",x"fb"),
  1223 => (x"87",x"ed",x"c1",x"05"),
  1224 => (x"4a",x"66",x"c0",x"c1"),
  1225 => (x"7e",x"6a",x"82",x"c4"),
  1226 => (x"dc",x"c1",x"1e",x"72"),
  1227 => (x"66",x"c4",x"48",x"f7"),
  1228 => (x"4a",x"a1",x"c8",x"49"),
  1229 => (x"aa",x"71",x"41",x"20"),
  1230 => (x"10",x"87",x"f9",x"05"),
  1231 => (x"c1",x"4a",x"26",x"51"),
  1232 => (x"c1",x"48",x"66",x"c0"),
  1233 => (x"6a",x"78",x"ee",x"c4"),
  1234 => (x"74",x"81",x"c7",x"49"),
  1235 => (x"66",x"c0",x"c1",x"51"),
  1236 => (x"c1",x"81",x"c8",x"49"),
  1237 => (x"66",x"c0",x"c1",x"51"),
  1238 => (x"c0",x"81",x"c9",x"49"),
  1239 => (x"66",x"c0",x"c1",x"51"),
  1240 => (x"c0",x"81",x"ca",x"49"),
  1241 => (x"d8",x"1e",x"c1",x"51"),
  1242 => (x"c8",x"49",x"6a",x"1e"),
  1243 => (x"87",x"c2",x"e3",x"81"),
  1244 => (x"c4",x"c1",x"86",x"c8"),
  1245 => (x"a8",x"c0",x"48",x"66"),
  1246 => (x"c8",x"87",x"c7",x"01"),
  1247 => (x"78",x"c1",x"48",x"a6"),
  1248 => (x"c4",x"c1",x"87",x"ce"),
  1249 => (x"88",x"c1",x"48",x"66"),
  1250 => (x"c3",x"58",x"a6",x"d0"),
  1251 => (x"87",x"ce",x"e2",x"87"),
  1252 => (x"c2",x"48",x"a6",x"d0"),
  1253 => (x"02",x"9c",x"74",x"78"),
  1254 => (x"c8",x"87",x"e3",x"cd"),
  1255 => (x"c8",x"c1",x"48",x"66"),
  1256 => (x"cd",x"03",x"a8",x"66"),
  1257 => (x"a6",x"dc",x"87",x"d8"),
  1258 => (x"e8",x"78",x"c0",x"48"),
  1259 => (x"e0",x"78",x"c0",x"80"),
  1260 => (x"4c",x"70",x"87",x"fc"),
  1261 => (x"05",x"ac",x"d0",x"c1"),
  1262 => (x"c4",x"87",x"d8",x"c2"),
  1263 => (x"e0",x"e3",x"7e",x"66"),
  1264 => (x"c8",x"49",x"70",x"87"),
  1265 => (x"e5",x"e0",x"59",x"a6"),
  1266 => (x"c0",x"4c",x"70",x"87"),
  1267 => (x"c1",x"05",x"ac",x"ec"),
  1268 => (x"66",x"c8",x"87",x"ec"),
  1269 => (x"c1",x"91",x"cb",x"49"),
  1270 => (x"c4",x"81",x"66",x"c0"),
  1271 => (x"4d",x"6a",x"4a",x"a1"),
  1272 => (x"c4",x"4a",x"a1",x"c8"),
  1273 => (x"c5",x"c1",x"52",x"66"),
  1274 => (x"c1",x"e0",x"79",x"ef"),
  1275 => (x"9c",x"4c",x"70",x"87"),
  1276 => (x"c0",x"87",x"d9",x"02"),
  1277 => (x"d3",x"02",x"ac",x"fb"),
  1278 => (x"ff",x"55",x"74",x"87"),
  1279 => (x"70",x"87",x"ef",x"df"),
  1280 => (x"c7",x"02",x"9c",x"4c"),
  1281 => (x"ac",x"fb",x"c0",x"87"),
  1282 => (x"87",x"ed",x"ff",x"05"),
  1283 => (x"c2",x"55",x"e0",x"c0"),
  1284 => (x"97",x"c0",x"55",x"c1"),
  1285 => (x"49",x"66",x"d8",x"7d"),
  1286 => (x"db",x"05",x"a9",x"6e"),
  1287 => (x"48",x"66",x"c8",x"87"),
  1288 => (x"04",x"a8",x"66",x"cc"),
  1289 => (x"66",x"c8",x"87",x"ca"),
  1290 => (x"cc",x"80",x"c1",x"48"),
  1291 => (x"87",x"c8",x"58",x"a6"),
  1292 => (x"c1",x"48",x"66",x"cc"),
  1293 => (x"58",x"a6",x"d0",x"88"),
  1294 => (x"87",x"f2",x"de",x"ff"),
  1295 => (x"d0",x"c1",x"4c",x"70"),
  1296 => (x"87",x"c8",x"05",x"ac"),
  1297 => (x"c1",x"48",x"66",x"d4"),
  1298 => (x"58",x"a6",x"d8",x"80"),
  1299 => (x"02",x"ac",x"d0",x"c1"),
  1300 => (x"c0",x"87",x"e8",x"fd"),
  1301 => (x"d8",x"48",x"a6",x"e0"),
  1302 => (x"66",x"c4",x"78",x"66"),
  1303 => (x"66",x"e0",x"c0",x"48"),
  1304 => (x"eb",x"c9",x"05",x"a8"),
  1305 => (x"a6",x"e4",x"c0",x"87"),
  1306 => (x"74",x"78",x"c0",x"48"),
  1307 => (x"88",x"fb",x"c0",x"48"),
  1308 => (x"98",x"48",x"7e",x"70"),
  1309 => (x"87",x"ed",x"c9",x"02"),
  1310 => (x"70",x"88",x"cb",x"48"),
  1311 => (x"02",x"98",x"48",x"7e"),
  1312 => (x"48",x"87",x"cd",x"c1"),
  1313 => (x"7e",x"70",x"88",x"c9"),
  1314 => (x"c4",x"02",x"98",x"48"),
  1315 => (x"c4",x"48",x"87",x"c1"),
  1316 => (x"48",x"7e",x"70",x"88"),
  1317 => (x"87",x"ce",x"02",x"98"),
  1318 => (x"70",x"88",x"c1",x"48"),
  1319 => (x"02",x"98",x"48",x"7e"),
  1320 => (x"c8",x"87",x"ec",x"c3"),
  1321 => (x"a6",x"dc",x"87",x"e1"),
  1322 => (x"78",x"f0",x"c0",x"48"),
  1323 => (x"87",x"fe",x"dc",x"ff"),
  1324 => (x"ec",x"c0",x"4c",x"70"),
  1325 => (x"c4",x"c0",x"02",x"ac"),
  1326 => (x"a6",x"e0",x"c0",x"87"),
  1327 => (x"ac",x"ec",x"c0",x"5c"),
  1328 => (x"ff",x"87",x"cd",x"02"),
  1329 => (x"70",x"87",x"e7",x"dc"),
  1330 => (x"ac",x"ec",x"c0",x"4c"),
  1331 => (x"87",x"f3",x"ff",x"05"),
  1332 => (x"02",x"ac",x"ec",x"c0"),
  1333 => (x"ff",x"87",x"c4",x"c0"),
  1334 => (x"c0",x"87",x"d3",x"dc"),
  1335 => (x"d0",x"1e",x"ca",x"1e"),
  1336 => (x"91",x"cb",x"49",x"66"),
  1337 => (x"48",x"66",x"c8",x"c1"),
  1338 => (x"a6",x"cc",x"80",x"71"),
  1339 => (x"48",x"66",x"c8",x"58"),
  1340 => (x"a6",x"d0",x"80",x"c4"),
  1341 => (x"bf",x"66",x"cc",x"58"),
  1342 => (x"f5",x"dc",x"ff",x"49"),
  1343 => (x"de",x"1e",x"c1",x"87"),
  1344 => (x"bf",x"66",x"d4",x"1e"),
  1345 => (x"e9",x"dc",x"ff",x"49"),
  1346 => (x"70",x"86",x"d0",x"87"),
  1347 => (x"89",x"09",x"c0",x"49"),
  1348 => (x"59",x"a6",x"ec",x"c0"),
  1349 => (x"48",x"66",x"e8",x"c0"),
  1350 => (x"c0",x"06",x"a8",x"c0"),
  1351 => (x"e8",x"c0",x"87",x"ee"),
  1352 => (x"a8",x"dd",x"48",x"66"),
  1353 => (x"87",x"e4",x"c0",x"03"),
  1354 => (x"49",x"bf",x"66",x"c4"),
  1355 => (x"81",x"66",x"e8",x"c0"),
  1356 => (x"c0",x"51",x"e0",x"c0"),
  1357 => (x"c1",x"49",x"66",x"e8"),
  1358 => (x"bf",x"66",x"c4",x"81"),
  1359 => (x"51",x"c1",x"c2",x"81"),
  1360 => (x"49",x"66",x"e8",x"c0"),
  1361 => (x"66",x"c4",x"81",x"c2"),
  1362 => (x"51",x"c0",x"81",x"bf"),
  1363 => (x"c4",x"c1",x"48",x"6e"),
  1364 => (x"49",x"6e",x"78",x"ee"),
  1365 => (x"66",x"d0",x"81",x"c8"),
  1366 => (x"c9",x"49",x"6e",x"51"),
  1367 => (x"51",x"66",x"d4",x"81"),
  1368 => (x"81",x"ca",x"49",x"6e"),
  1369 => (x"d0",x"51",x"66",x"dc"),
  1370 => (x"80",x"c1",x"48",x"66"),
  1371 => (x"c8",x"58",x"a6",x"d4"),
  1372 => (x"66",x"cc",x"48",x"66"),
  1373 => (x"cb",x"c0",x"04",x"a8"),
  1374 => (x"48",x"66",x"c8",x"87"),
  1375 => (x"a6",x"cc",x"80",x"c1"),
  1376 => (x"87",x"e1",x"c5",x"58"),
  1377 => (x"c1",x"48",x"66",x"cc"),
  1378 => (x"58",x"a6",x"d0",x"88"),
  1379 => (x"ff",x"87",x"d6",x"c5"),
  1380 => (x"70",x"87",x"ce",x"dc"),
  1381 => (x"a6",x"ec",x"c0",x"49"),
  1382 => (x"c4",x"dc",x"ff",x"59"),
  1383 => (x"c0",x"49",x"70",x"87"),
  1384 => (x"dc",x"59",x"a6",x"e0"),
  1385 => (x"ec",x"c0",x"48",x"66"),
  1386 => (x"ca",x"c0",x"05",x"a8"),
  1387 => (x"48",x"a6",x"dc",x"87"),
  1388 => (x"78",x"66",x"e8",x"c0"),
  1389 => (x"ff",x"87",x"c4",x"c0"),
  1390 => (x"c8",x"87",x"f3",x"d8"),
  1391 => (x"91",x"cb",x"49",x"66"),
  1392 => (x"48",x"66",x"c0",x"c1"),
  1393 => (x"7e",x"70",x"80",x"71"),
  1394 => (x"6e",x"82",x"c8",x"4a"),
  1395 => (x"c0",x"81",x"ca",x"49"),
  1396 => (x"dc",x"51",x"66",x"e8"),
  1397 => (x"81",x"c1",x"49",x"66"),
  1398 => (x"89",x"66",x"e8",x"c0"),
  1399 => (x"30",x"71",x"48",x"c1"),
  1400 => (x"89",x"c1",x"49",x"70"),
  1401 => (x"c2",x"7a",x"97",x"71"),
  1402 => (x"49",x"bf",x"e8",x"f3"),
  1403 => (x"29",x"66",x"e8",x"c0"),
  1404 => (x"48",x"4a",x"6a",x"97"),
  1405 => (x"f0",x"c0",x"98",x"71"),
  1406 => (x"49",x"6e",x"58",x"a6"),
  1407 => (x"4d",x"69",x"81",x"c4"),
  1408 => (x"48",x"66",x"e0",x"c0"),
  1409 => (x"02",x"a8",x"66",x"c4"),
  1410 => (x"c4",x"87",x"c8",x"c0"),
  1411 => (x"78",x"c0",x"48",x"a6"),
  1412 => (x"c4",x"87",x"c5",x"c0"),
  1413 => (x"78",x"c1",x"48",x"a6"),
  1414 => (x"c0",x"1e",x"66",x"c4"),
  1415 => (x"49",x"75",x"1e",x"e0"),
  1416 => (x"87",x"ce",x"d8",x"ff"),
  1417 => (x"4c",x"70",x"86",x"c8"),
  1418 => (x"06",x"ac",x"b7",x"c0"),
  1419 => (x"74",x"87",x"d4",x"c1"),
  1420 => (x"49",x"e0",x"c0",x"85"),
  1421 => (x"4b",x"75",x"89",x"74"),
  1422 => (x"4a",x"c0",x"dd",x"c1"),
  1423 => (x"e6",x"e9",x"fe",x"71"),
  1424 => (x"c0",x"85",x"c2",x"87"),
  1425 => (x"c1",x"48",x"66",x"e4"),
  1426 => (x"a6",x"e8",x"c0",x"80"),
  1427 => (x"66",x"ec",x"c0",x"58"),
  1428 => (x"70",x"81",x"c1",x"49"),
  1429 => (x"c8",x"c0",x"02",x"a9"),
  1430 => (x"48",x"a6",x"c4",x"87"),
  1431 => (x"c5",x"c0",x"78",x"c0"),
  1432 => (x"48",x"a6",x"c4",x"87"),
  1433 => (x"66",x"c4",x"78",x"c1"),
  1434 => (x"49",x"a4",x"c2",x"1e"),
  1435 => (x"71",x"48",x"e0",x"c0"),
  1436 => (x"1e",x"49",x"70",x"88"),
  1437 => (x"d6",x"ff",x"49",x"75"),
  1438 => (x"86",x"c8",x"87",x"f8"),
  1439 => (x"01",x"a8",x"b7",x"c0"),
  1440 => (x"c0",x"87",x"c0",x"ff"),
  1441 => (x"c0",x"02",x"66",x"e4"),
  1442 => (x"49",x"6e",x"87",x"d1"),
  1443 => (x"e4",x"c0",x"81",x"c9"),
  1444 => (x"48",x"6e",x"51",x"66"),
  1445 => (x"78",x"ff",x"c6",x"c1"),
  1446 => (x"6e",x"87",x"cc",x"c0"),
  1447 => (x"c2",x"81",x"c9",x"49"),
  1448 => (x"c1",x"48",x"6e",x"51"),
  1449 => (x"c8",x"78",x"ee",x"c8"),
  1450 => (x"66",x"cc",x"48",x"66"),
  1451 => (x"cb",x"c0",x"04",x"a8"),
  1452 => (x"48",x"66",x"c8",x"87"),
  1453 => (x"a6",x"cc",x"80",x"c1"),
  1454 => (x"87",x"e9",x"c0",x"58"),
  1455 => (x"c1",x"48",x"66",x"cc"),
  1456 => (x"58",x"a6",x"d0",x"88"),
  1457 => (x"ff",x"87",x"de",x"c0"),
  1458 => (x"70",x"87",x"d3",x"d5"),
  1459 => (x"87",x"d5",x"c0",x"4c"),
  1460 => (x"05",x"ac",x"c6",x"c1"),
  1461 => (x"d0",x"87",x"c8",x"c0"),
  1462 => (x"80",x"c1",x"48",x"66"),
  1463 => (x"ff",x"58",x"a6",x"d4"),
  1464 => (x"70",x"87",x"fb",x"d4"),
  1465 => (x"48",x"66",x"d4",x"4c"),
  1466 => (x"a6",x"d8",x"80",x"c1"),
  1467 => (x"02",x"9c",x"74",x"58"),
  1468 => (x"c8",x"87",x"cb",x"c0"),
  1469 => (x"c8",x"c1",x"48",x"66"),
  1470 => (x"f2",x"04",x"a8",x"66"),
  1471 => (x"d4",x"ff",x"87",x"e8"),
  1472 => (x"66",x"c8",x"87",x"d3"),
  1473 => (x"03",x"a8",x"c7",x"48"),
  1474 => (x"c2",x"87",x"e5",x"c0"),
  1475 => (x"c0",x"48",x"fc",x"ef"),
  1476 => (x"49",x"66",x"c8",x"78"),
  1477 => (x"c0",x"c1",x"91",x"cb"),
  1478 => (x"a1",x"c4",x"81",x"66"),
  1479 => (x"c0",x"4a",x"6a",x"4a"),
  1480 => (x"66",x"c8",x"79",x"52"),
  1481 => (x"cc",x"80",x"c1",x"48"),
  1482 => (x"a8",x"c7",x"58",x"a6"),
  1483 => (x"87",x"db",x"ff",x"04"),
  1484 => (x"ff",x"8e",x"d0",x"ff"),
  1485 => (x"4c",x"87",x"e5",x"de"),
  1486 => (x"20",x"64",x"61",x"6f"),
  1487 => (x"00",x"20",x"2e",x"2a"),
  1488 => (x"1e",x"00",x"20",x"3a"),
  1489 => (x"4b",x"71",x"1e",x"73"),
  1490 => (x"87",x"c6",x"02",x"9b"),
  1491 => (x"48",x"f8",x"ef",x"c2"),
  1492 => (x"1e",x"c7",x"78",x"c0"),
  1493 => (x"bf",x"f8",x"ef",x"c2"),
  1494 => (x"e1",x"c1",x"1e",x"49"),
  1495 => (x"ef",x"c2",x"1e",x"d0"),
  1496 => (x"ed",x"49",x"bf",x"e0"),
  1497 => (x"86",x"cc",x"87",x"e8"),
  1498 => (x"bf",x"e0",x"ef",x"c2"),
  1499 => (x"87",x"e7",x"e8",x"49"),
  1500 => (x"c8",x"02",x"9b",x"73"),
  1501 => (x"d0",x"e1",x"c1",x"87"),
  1502 => (x"c6",x"e3",x"c0",x"49"),
  1503 => (x"df",x"dd",x"ff",x"87"),
  1504 => (x"1e",x"73",x"1e",x"87"),
  1505 => (x"e0",x"c1",x"4b",x"c0"),
  1506 => (x"50",x"c0",x"48",x"fc"),
  1507 => (x"bf",x"f3",x"e2",x"c1"),
  1508 => (x"d9",x"d8",x"ff",x"49"),
  1509 => (x"05",x"98",x"70",x"87"),
  1510 => (x"de",x"c1",x"87",x"c4"),
  1511 => (x"48",x"73",x"4b",x"e4"),
  1512 => (x"87",x"fc",x"dc",x"ff"),
  1513 => (x"20",x"4d",x"4f",x"52"),
  1514 => (x"64",x"61",x"6f",x"6c"),
  1515 => (x"20",x"67",x"6e",x"69"),
  1516 => (x"6c",x"69",x"61",x"66"),
  1517 => (x"1e",x"00",x"64",x"65"),
  1518 => (x"c1",x"87",x"df",x"c7"),
  1519 => (x"87",x"c3",x"fe",x"49"),
  1520 => (x"87",x"c9",x"ed",x"fe"),
  1521 => (x"cd",x"02",x"98",x"70"),
  1522 => (x"e2",x"f4",x"fe",x"87"),
  1523 => (x"02",x"98",x"70",x"87"),
  1524 => (x"4a",x"c1",x"87",x"c4"),
  1525 => (x"4a",x"c0",x"87",x"c2"),
  1526 => (x"ce",x"05",x"9a",x"72"),
  1527 => (x"c1",x"1e",x"c0",x"87"),
  1528 => (x"c0",x"49",x"c7",x"e0"),
  1529 => (x"c4",x"87",x"d3",x"ee"),
  1530 => (x"c0",x"87",x"fe",x"86"),
  1531 => (x"d2",x"e0",x"c1",x"1e"),
  1532 => (x"c5",x"ee",x"c0",x"49"),
  1533 => (x"fe",x"1e",x"c0",x"87"),
  1534 => (x"49",x"70",x"87",x"c7"),
  1535 => (x"87",x"fa",x"ed",x"c0"),
  1536 => (x"f8",x"87",x"d6",x"c3"),
  1537 => (x"53",x"4f",x"26",x"8e"),
  1538 => (x"61",x"66",x"20",x"44"),
  1539 => (x"64",x"65",x"6c",x"69"),
  1540 => (x"6f",x"42",x"00",x"2e"),
  1541 => (x"6e",x"69",x"74",x"6f"),
  1542 => (x"2e",x"2e",x"2e",x"67"),
  1543 => (x"e5",x"c0",x"1e",x"00"),
  1544 => (x"87",x"fa",x"87",x"df"),
  1545 => (x"c2",x"1e",x"4f",x"26"),
  1546 => (x"c0",x"48",x"f8",x"ef"),
  1547 => (x"e0",x"ef",x"c2",x"78"),
  1548 => (x"fe",x"78",x"c0",x"48"),
  1549 => (x"87",x"e5",x"87",x"c1"),
  1550 => (x"4f",x"26",x"48",x"c0"),
  1551 => (x"00",x"01",x"00",x"00"),
  1552 => (x"20",x"80",x"00",x"00"),
  1553 => (x"74",x"69",x"78",x"45"),
  1554 => (x"42",x"20",x"80",x"00"),
  1555 => (x"00",x"6b",x"63",x"61"),
  1556 => (x"00",x"00",x"0f",x"32"),
  1557 => (x"00",x"00",x"2c",x"0c"),
  1558 => (x"32",x"00",x"00",x"00"),
  1559 => (x"2a",x"00",x"00",x"0f"),
  1560 => (x"00",x"00",x"00",x"2c"),
  1561 => (x"0f",x"32",x"00",x"00"),
  1562 => (x"2c",x"48",x"00",x"00"),
  1563 => (x"00",x"00",x"00",x"00"),
  1564 => (x"00",x"0f",x"32",x"00"),
  1565 => (x"00",x"2c",x"66",x"00"),
  1566 => (x"00",x"00",x"00",x"00"),
  1567 => (x"00",x"00",x"0f",x"32"),
  1568 => (x"00",x"00",x"2c",x"84"),
  1569 => (x"32",x"00",x"00",x"00"),
  1570 => (x"a2",x"00",x"00",x"0f"),
  1571 => (x"00",x"00",x"00",x"2c"),
  1572 => (x"0f",x"32",x"00",x"00"),
  1573 => (x"2c",x"c0",x"00",x"00"),
  1574 => (x"00",x"00",x"00",x"00"),
  1575 => (x"00",x"11",x"6f",x"00"),
  1576 => (x"00",x"00",x"00",x"00"),
  1577 => (x"00",x"00",x"00",x"00"),
  1578 => (x"00",x"00",x"12",x"3f"),
  1579 => (x"00",x"00",x"00",x"00"),
  1580 => (x"b7",x"00",x"00",x"00"),
  1581 => (x"50",x"00",x"00",x"18"),
  1582 => (x"30",x"32",x"54",x"45"),
  1583 => (x"52",x"20",x"31",x"30"),
  1584 => (x"1e",x"00",x"4d",x"4f"),
  1585 => (x"c0",x"48",x"f0",x"fe"),
  1586 => (x"79",x"09",x"cd",x"78"),
  1587 => (x"1e",x"4f",x"26",x"09"),
  1588 => (x"bf",x"f0",x"fe",x"1e"),
  1589 => (x"26",x"26",x"48",x"7e"),
  1590 => (x"f0",x"fe",x"1e",x"4f"),
  1591 => (x"26",x"78",x"c1",x"48"),
  1592 => (x"f0",x"fe",x"1e",x"4f"),
  1593 => (x"26",x"78",x"c0",x"48"),
  1594 => (x"4a",x"71",x"1e",x"4f"),
  1595 => (x"26",x"52",x"52",x"c0"),
  1596 => (x"5b",x"5e",x"0e",x"4f"),
  1597 => (x"f4",x"0e",x"5d",x"5c"),
  1598 => (x"97",x"4d",x"71",x"86"),
  1599 => (x"a5",x"c1",x"7e",x"6d"),
  1600 => (x"48",x"6c",x"97",x"4c"),
  1601 => (x"6e",x"58",x"a6",x"c8"),
  1602 => (x"a8",x"66",x"c4",x"48"),
  1603 => (x"ff",x"87",x"c5",x"05"),
  1604 => (x"87",x"e6",x"c0",x"48"),
  1605 => (x"c2",x"87",x"ca",x"ff"),
  1606 => (x"6c",x"97",x"49",x"a5"),
  1607 => (x"4b",x"a3",x"71",x"4b"),
  1608 => (x"97",x"4b",x"6b",x"97"),
  1609 => (x"48",x"6e",x"7e",x"6c"),
  1610 => (x"a6",x"c8",x"80",x"c1"),
  1611 => (x"cc",x"98",x"c7",x"58"),
  1612 => (x"97",x"70",x"58",x"a6"),
  1613 => (x"87",x"e1",x"fe",x"7c"),
  1614 => (x"8e",x"f4",x"48",x"73"),
  1615 => (x"4c",x"26",x"4d",x"26"),
  1616 => (x"4f",x"26",x"4b",x"26"),
  1617 => (x"5c",x"5b",x"5e",x"0e"),
  1618 => (x"71",x"86",x"f4",x"0e"),
  1619 => (x"4a",x"66",x"d8",x"4c"),
  1620 => (x"c2",x"9a",x"ff",x"c3"),
  1621 => (x"6c",x"97",x"4b",x"a4"),
  1622 => (x"49",x"a1",x"73",x"49"),
  1623 => (x"6c",x"97",x"51",x"72"),
  1624 => (x"c1",x"48",x"6e",x"7e"),
  1625 => (x"58",x"a6",x"c8",x"80"),
  1626 => (x"a6",x"cc",x"98",x"c7"),
  1627 => (x"f4",x"54",x"70",x"58"),
  1628 => (x"87",x"ca",x"ff",x"8e"),
  1629 => (x"e8",x"fd",x"1e",x"1e"),
  1630 => (x"4a",x"bf",x"e0",x"87"),
  1631 => (x"c0",x"e0",x"c0",x"49"),
  1632 => (x"87",x"cb",x"02",x"99"),
  1633 => (x"f3",x"c2",x"1e",x"72"),
  1634 => (x"f7",x"fe",x"49",x"de"),
  1635 => (x"fc",x"86",x"c4",x"87"),
  1636 => (x"7e",x"70",x"87",x"fd"),
  1637 => (x"26",x"87",x"c2",x"fd"),
  1638 => (x"c2",x"1e",x"4f",x"26"),
  1639 => (x"fd",x"49",x"de",x"f3"),
  1640 => (x"e5",x"c1",x"87",x"c7"),
  1641 => (x"da",x"fc",x"49",x"f4"),
  1642 => (x"87",x"ee",x"c3",x"87"),
  1643 => (x"5e",x"0e",x"4f",x"26"),
  1644 => (x"0e",x"5d",x"5c",x"5b"),
  1645 => (x"f3",x"c2",x"4d",x"71"),
  1646 => (x"f4",x"fc",x"49",x"de"),
  1647 => (x"c0",x"4b",x"70",x"87"),
  1648 => (x"c3",x"04",x"ab",x"b7"),
  1649 => (x"f0",x"c3",x"87",x"c2"),
  1650 => (x"87",x"c9",x"05",x"ab"),
  1651 => (x"48",x"d2",x"ea",x"c1"),
  1652 => (x"e3",x"c2",x"78",x"c1"),
  1653 => (x"ab",x"e0",x"c3",x"87"),
  1654 => (x"c1",x"87",x"c9",x"05"),
  1655 => (x"c1",x"48",x"d6",x"ea"),
  1656 => (x"87",x"d4",x"c2",x"78"),
  1657 => (x"bf",x"d6",x"ea",x"c1"),
  1658 => (x"c2",x"87",x"c6",x"02"),
  1659 => (x"c2",x"4c",x"a3",x"c0"),
  1660 => (x"c1",x"4c",x"73",x"87"),
  1661 => (x"02",x"bf",x"d2",x"ea"),
  1662 => (x"74",x"87",x"e0",x"c0"),
  1663 => (x"29",x"b7",x"c4",x"49"),
  1664 => (x"e9",x"eb",x"c1",x"91"),
  1665 => (x"cf",x"4a",x"74",x"81"),
  1666 => (x"c1",x"92",x"c2",x"9a"),
  1667 => (x"70",x"30",x"72",x"48"),
  1668 => (x"72",x"ba",x"ff",x"4a"),
  1669 => (x"70",x"98",x"69",x"48"),
  1670 => (x"74",x"87",x"db",x"79"),
  1671 => (x"29",x"b7",x"c4",x"49"),
  1672 => (x"e9",x"eb",x"c1",x"91"),
  1673 => (x"cf",x"4a",x"74",x"81"),
  1674 => (x"c3",x"92",x"c2",x"9a"),
  1675 => (x"70",x"30",x"72",x"48"),
  1676 => (x"b0",x"69",x"48",x"4a"),
  1677 => (x"9d",x"75",x"79",x"70"),
  1678 => (x"87",x"f0",x"c0",x"05"),
  1679 => (x"c8",x"48",x"d0",x"ff"),
  1680 => (x"d4",x"ff",x"78",x"e1"),
  1681 => (x"c1",x"78",x"c5",x"48"),
  1682 => (x"02",x"bf",x"d6",x"ea"),
  1683 => (x"e0",x"c3",x"87",x"c3"),
  1684 => (x"d2",x"ea",x"c1",x"78"),
  1685 => (x"87",x"c6",x"02",x"bf"),
  1686 => (x"c3",x"48",x"d4",x"ff"),
  1687 => (x"d4",x"ff",x"78",x"f0"),
  1688 => (x"ff",x"78",x"73",x"48"),
  1689 => (x"e1",x"c8",x"48",x"d0"),
  1690 => (x"78",x"e0",x"c0",x"78"),
  1691 => (x"48",x"d6",x"ea",x"c1"),
  1692 => (x"ea",x"c1",x"78",x"c0"),
  1693 => (x"78",x"c0",x"48",x"d2"),
  1694 => (x"49",x"de",x"f3",x"c2"),
  1695 => (x"70",x"87",x"f2",x"f9"),
  1696 => (x"ab",x"b7",x"c0",x"4b"),
  1697 => (x"87",x"fe",x"fc",x"03"),
  1698 => (x"4d",x"26",x"48",x"c0"),
  1699 => (x"4b",x"26",x"4c",x"26"),
  1700 => (x"00",x"00",x"4f",x"26"),
  1701 => (x"00",x"00",x"00",x"00"),
  1702 => (x"c0",x"1e",x"00",x"00"),
  1703 => (x"c4",x"49",x"72",x"4a"),
  1704 => (x"e9",x"eb",x"c1",x"91"),
  1705 => (x"c1",x"79",x"c0",x"81"),
  1706 => (x"aa",x"b7",x"d0",x"82"),
  1707 => (x"26",x"87",x"ee",x"04"),
  1708 => (x"5b",x"5e",x"0e",x"4f"),
  1709 => (x"71",x"0e",x"5d",x"5c"),
  1710 => (x"87",x"e5",x"f8",x"4d"),
  1711 => (x"b7",x"c4",x"4a",x"75"),
  1712 => (x"eb",x"c1",x"92",x"2a"),
  1713 => (x"4c",x"75",x"82",x"e9"),
  1714 => (x"94",x"c2",x"9c",x"cf"),
  1715 => (x"74",x"4b",x"49",x"6a"),
  1716 => (x"c2",x"9b",x"c3",x"2b"),
  1717 => (x"70",x"30",x"74",x"48"),
  1718 => (x"74",x"bc",x"ff",x"4c"),
  1719 => (x"70",x"98",x"71",x"48"),
  1720 => (x"87",x"f5",x"f7",x"7a"),
  1721 => (x"e1",x"fe",x"48",x"73"),
  1722 => (x"00",x"00",x"00",x"87"),
  1723 => (x"00",x"00",x"00",x"00"),
  1724 => (x"00",x"00",x"00",x"00"),
  1725 => (x"00",x"00",x"00",x"00"),
  1726 => (x"00",x"00",x"00",x"00"),
  1727 => (x"00",x"00",x"00",x"00"),
  1728 => (x"00",x"00",x"00",x"00"),
  1729 => (x"00",x"00",x"00",x"00"),
  1730 => (x"00",x"00",x"00",x"00"),
  1731 => (x"00",x"00",x"00",x"00"),
  1732 => (x"00",x"00",x"00",x"00"),
  1733 => (x"00",x"00",x"00",x"00"),
  1734 => (x"00",x"00",x"00",x"00"),
  1735 => (x"00",x"00",x"00",x"00"),
  1736 => (x"00",x"00",x"00",x"00"),
  1737 => (x"00",x"00",x"00",x"00"),
  1738 => (x"d0",x"ff",x"1e",x"00"),
  1739 => (x"78",x"e1",x"c8",x"48"),
  1740 => (x"d4",x"ff",x"48",x"71"),
  1741 => (x"66",x"c4",x"78",x"08"),
  1742 => (x"08",x"d4",x"ff",x"48"),
  1743 => (x"1e",x"4f",x"26",x"78"),
  1744 => (x"66",x"c4",x"4a",x"71"),
  1745 => (x"49",x"72",x"1e",x"49"),
  1746 => (x"ff",x"87",x"de",x"ff"),
  1747 => (x"e0",x"c0",x"48",x"d0"),
  1748 => (x"4f",x"26",x"26",x"78"),
  1749 => (x"71",x"1e",x"73",x"1e"),
  1750 => (x"49",x"66",x"c8",x"4b"),
  1751 => (x"c1",x"4a",x"73",x"1e"),
  1752 => (x"ff",x"49",x"a2",x"e0"),
  1753 => (x"c4",x"26",x"87",x"d9"),
  1754 => (x"26",x"4d",x"26",x"87"),
  1755 => (x"26",x"4b",x"26",x"4c"),
  1756 => (x"d4",x"ff",x"1e",x"4f"),
  1757 => (x"7a",x"ff",x"c3",x"4a"),
  1758 => (x"c0",x"48",x"d0",x"ff"),
  1759 => (x"7a",x"de",x"78",x"e1"),
  1760 => (x"bf",x"e8",x"f3",x"c2"),
  1761 => (x"c8",x"48",x"49",x"7a"),
  1762 => (x"71",x"7a",x"70",x"28"),
  1763 => (x"70",x"28",x"d0",x"48"),
  1764 => (x"d8",x"48",x"71",x"7a"),
  1765 => (x"ff",x"7a",x"70",x"28"),
  1766 => (x"e0",x"c0",x"48",x"d0"),
  1767 => (x"1e",x"4f",x"26",x"78"),
  1768 => (x"c8",x"48",x"d0",x"ff"),
  1769 => (x"48",x"71",x"78",x"c9"),
  1770 => (x"78",x"08",x"d4",x"ff"),
  1771 => (x"71",x"1e",x"4f",x"26"),
  1772 => (x"87",x"eb",x"49",x"4a"),
  1773 => (x"c8",x"48",x"d0",x"ff"),
  1774 => (x"1e",x"4f",x"26",x"78"),
  1775 => (x"4b",x"71",x"1e",x"73"),
  1776 => (x"bf",x"f8",x"f3",x"c2"),
  1777 => (x"c2",x"87",x"c3",x"02"),
  1778 => (x"d0",x"ff",x"87",x"eb"),
  1779 => (x"78",x"c9",x"c8",x"48"),
  1780 => (x"e0",x"c0",x"49",x"73"),
  1781 => (x"48",x"d4",x"ff",x"b1"),
  1782 => (x"f3",x"c2",x"78",x"71"),
  1783 => (x"78",x"c0",x"48",x"ec"),
  1784 => (x"c5",x"02",x"66",x"c8"),
  1785 => (x"49",x"ff",x"c3",x"87"),
  1786 => (x"49",x"c0",x"87",x"c2"),
  1787 => (x"59",x"f4",x"f3",x"c2"),
  1788 => (x"c6",x"02",x"66",x"cc"),
  1789 => (x"d5",x"d5",x"c5",x"87"),
  1790 => (x"cf",x"87",x"c4",x"4a"),
  1791 => (x"c2",x"4a",x"ff",x"ff"),
  1792 => (x"c2",x"5a",x"f8",x"f3"),
  1793 => (x"c1",x"48",x"f8",x"f3"),
  1794 => (x"26",x"87",x"c4",x"78"),
  1795 => (x"26",x"4c",x"26",x"4d"),
  1796 => (x"0e",x"4f",x"26",x"4b"),
  1797 => (x"5d",x"5c",x"5b",x"5e"),
  1798 => (x"c2",x"4a",x"71",x"0e"),
  1799 => (x"4c",x"bf",x"f4",x"f3"),
  1800 => (x"cb",x"02",x"9a",x"72"),
  1801 => (x"91",x"c8",x"49",x"87"),
  1802 => (x"4b",x"f1",x"ee",x"c1"),
  1803 => (x"87",x"c4",x"83",x"71"),
  1804 => (x"4b",x"f1",x"f2",x"c1"),
  1805 => (x"49",x"13",x"4d",x"c0"),
  1806 => (x"f3",x"c2",x"99",x"74"),
  1807 => (x"ff",x"b9",x"bf",x"f0"),
  1808 => (x"78",x"71",x"48",x"d4"),
  1809 => (x"85",x"2c",x"b7",x"c1"),
  1810 => (x"04",x"ad",x"b7",x"c8"),
  1811 => (x"f3",x"c2",x"87",x"e8"),
  1812 => (x"c8",x"48",x"bf",x"ec"),
  1813 => (x"f0",x"f3",x"c2",x"80"),
  1814 => (x"87",x"ef",x"fe",x"58"),
  1815 => (x"71",x"1e",x"73",x"1e"),
  1816 => (x"9a",x"4a",x"13",x"4b"),
  1817 => (x"72",x"87",x"cb",x"02"),
  1818 => (x"87",x"e7",x"fe",x"49"),
  1819 => (x"05",x"9a",x"4a",x"13"),
  1820 => (x"da",x"fe",x"87",x"f5"),
  1821 => (x"f3",x"c2",x"1e",x"87"),
  1822 => (x"c2",x"49",x"bf",x"ec"),
  1823 => (x"c1",x"48",x"ec",x"f3"),
  1824 => (x"c0",x"c4",x"78",x"a1"),
  1825 => (x"db",x"03",x"a9",x"b7"),
  1826 => (x"48",x"d4",x"ff",x"87"),
  1827 => (x"bf",x"f0",x"f3",x"c2"),
  1828 => (x"ec",x"f3",x"c2",x"78"),
  1829 => (x"f3",x"c2",x"49",x"bf"),
  1830 => (x"a1",x"c1",x"48",x"ec"),
  1831 => (x"b7",x"c0",x"c4",x"78"),
  1832 => (x"87",x"e5",x"04",x"a9"),
  1833 => (x"c8",x"48",x"d0",x"ff"),
  1834 => (x"f8",x"f3",x"c2",x"78"),
  1835 => (x"26",x"78",x"c0",x"48"),
  1836 => (x"00",x"00",x"00",x"4f"),
  1837 => (x"00",x"00",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"00",x"00",x"5f",x"5f"),
  1840 => (x"03",x"03",x"00",x"00"),
  1841 => (x"00",x"03",x"03",x"00"),
  1842 => (x"7f",x"7f",x"14",x"00"),
  1843 => (x"14",x"7f",x"7f",x"14"),
  1844 => (x"2e",x"24",x"00",x"00"),
  1845 => (x"12",x"3a",x"6b",x"6b"),
  1846 => (x"36",x"6a",x"4c",x"00"),
  1847 => (x"32",x"56",x"6c",x"18"),
  1848 => (x"4f",x"7e",x"30",x"00"),
  1849 => (x"68",x"3a",x"77",x"59"),
  1850 => (x"04",x"00",x"00",x"40"),
  1851 => (x"00",x"00",x"03",x"07"),
  1852 => (x"1c",x"00",x"00",x"00"),
  1853 => (x"00",x"41",x"63",x"3e"),
  1854 => (x"41",x"00",x"00",x"00"),
  1855 => (x"00",x"1c",x"3e",x"63"),
  1856 => (x"3e",x"2a",x"08",x"00"),
  1857 => (x"2a",x"3e",x"1c",x"1c"),
  1858 => (x"08",x"08",x"00",x"08"),
  1859 => (x"08",x"08",x"3e",x"3e"),
  1860 => (x"80",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"60",x"e0"),
  1862 => (x"08",x"08",x"00",x"00"),
  1863 => (x"08",x"08",x"08",x"08"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"60",x"60"),
  1866 => (x"30",x"60",x"40",x"00"),
  1867 => (x"03",x"06",x"0c",x"18"),
  1868 => (x"7f",x"3e",x"00",x"01"),
  1869 => (x"3e",x"7f",x"4d",x"59"),
  1870 => (x"06",x"04",x"00",x"00"),
  1871 => (x"00",x"00",x"7f",x"7f"),
  1872 => (x"63",x"42",x"00",x"00"),
  1873 => (x"46",x"4f",x"59",x"71"),
  1874 => (x"63",x"22",x"00",x"00"),
  1875 => (x"36",x"7f",x"49",x"49"),
  1876 => (x"16",x"1c",x"18",x"00"),
  1877 => (x"10",x"7f",x"7f",x"13"),
  1878 => (x"67",x"27",x"00",x"00"),
  1879 => (x"39",x"7d",x"45",x"45"),
  1880 => (x"7e",x"3c",x"00",x"00"),
  1881 => (x"30",x"79",x"49",x"4b"),
  1882 => (x"01",x"01",x"00",x"00"),
  1883 => (x"07",x"0f",x"79",x"71"),
  1884 => (x"7f",x"36",x"00",x"00"),
  1885 => (x"36",x"7f",x"49",x"49"),
  1886 => (x"4f",x"06",x"00",x"00"),
  1887 => (x"1e",x"3f",x"69",x"49"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"66",x"66"),
  1890 => (x"80",x"00",x"00",x"00"),
  1891 => (x"00",x"00",x"66",x"e6"),
  1892 => (x"08",x"08",x"00",x"00"),
  1893 => (x"22",x"22",x"14",x"14"),
  1894 => (x"14",x"14",x"00",x"00"),
  1895 => (x"14",x"14",x"14",x"14"),
  1896 => (x"22",x"22",x"00",x"00"),
  1897 => (x"08",x"08",x"14",x"14"),
  1898 => (x"03",x"02",x"00",x"00"),
  1899 => (x"06",x"0f",x"59",x"51"),
  1900 => (x"41",x"7f",x"3e",x"00"),
  1901 => (x"1e",x"1f",x"55",x"5d"),
  1902 => (x"7f",x"7e",x"00",x"00"),
  1903 => (x"7e",x"7f",x"09",x"09"),
  1904 => (x"7f",x"7f",x"00",x"00"),
  1905 => (x"36",x"7f",x"49",x"49"),
  1906 => (x"3e",x"1c",x"00",x"00"),
  1907 => (x"41",x"41",x"41",x"63"),
  1908 => (x"7f",x"7f",x"00",x"00"),
  1909 => (x"1c",x"3e",x"63",x"41"),
  1910 => (x"7f",x"7f",x"00",x"00"),
  1911 => (x"41",x"41",x"49",x"49"),
  1912 => (x"7f",x"7f",x"00",x"00"),
  1913 => (x"01",x"01",x"09",x"09"),
  1914 => (x"7f",x"3e",x"00",x"00"),
  1915 => (x"7a",x"7b",x"49",x"41"),
  1916 => (x"7f",x"7f",x"00",x"00"),
  1917 => (x"7f",x"7f",x"08",x"08"),
  1918 => (x"41",x"00",x"00",x"00"),
  1919 => (x"00",x"41",x"7f",x"7f"),
  1920 => (x"60",x"20",x"00",x"00"),
  1921 => (x"3f",x"7f",x"40",x"40"),
  1922 => (x"08",x"7f",x"7f",x"00"),
  1923 => (x"41",x"63",x"36",x"1c"),
  1924 => (x"7f",x"7f",x"00",x"00"),
  1925 => (x"40",x"40",x"40",x"40"),
  1926 => (x"06",x"7f",x"7f",x"00"),
  1927 => (x"7f",x"7f",x"06",x"0c"),
  1928 => (x"06",x"7f",x"7f",x"00"),
  1929 => (x"7f",x"7f",x"18",x"0c"),
  1930 => (x"7f",x"3e",x"00",x"00"),
  1931 => (x"3e",x"7f",x"41",x"41"),
  1932 => (x"7f",x"7f",x"00",x"00"),
  1933 => (x"06",x"0f",x"09",x"09"),
  1934 => (x"41",x"7f",x"3e",x"00"),
  1935 => (x"40",x"7e",x"7f",x"61"),
  1936 => (x"7f",x"7f",x"00",x"00"),
  1937 => (x"66",x"7f",x"19",x"09"),
  1938 => (x"6f",x"26",x"00",x"00"),
  1939 => (x"32",x"7b",x"59",x"4d"),
  1940 => (x"01",x"01",x"00",x"00"),
  1941 => (x"01",x"01",x"7f",x"7f"),
  1942 => (x"7f",x"3f",x"00",x"00"),
  1943 => (x"3f",x"7f",x"40",x"40"),
  1944 => (x"3f",x"0f",x"00",x"00"),
  1945 => (x"0f",x"3f",x"70",x"70"),
  1946 => (x"30",x"7f",x"7f",x"00"),
  1947 => (x"7f",x"7f",x"30",x"18"),
  1948 => (x"36",x"63",x"41",x"00"),
  1949 => (x"63",x"36",x"1c",x"1c"),
  1950 => (x"06",x"03",x"01",x"41"),
  1951 => (x"03",x"06",x"7c",x"7c"),
  1952 => (x"59",x"71",x"61",x"01"),
  1953 => (x"41",x"43",x"47",x"4d"),
  1954 => (x"7f",x"00",x"00",x"00"),
  1955 => (x"00",x"41",x"41",x"7f"),
  1956 => (x"06",x"03",x"01",x"00"),
  1957 => (x"60",x"30",x"18",x"0c"),
  1958 => (x"41",x"00",x"00",x"40"),
  1959 => (x"00",x"7f",x"7f",x"41"),
  1960 => (x"06",x"0c",x"08",x"00"),
  1961 => (x"08",x"0c",x"06",x"03"),
  1962 => (x"80",x"80",x"80",x"00"),
  1963 => (x"80",x"80",x"80",x"80"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"00",x"04",x"07",x"03"),
  1966 => (x"74",x"20",x"00",x"00"),
  1967 => (x"78",x"7c",x"54",x"54"),
  1968 => (x"7f",x"7f",x"00",x"00"),
  1969 => (x"38",x"7c",x"44",x"44"),
  1970 => (x"7c",x"38",x"00",x"00"),
  1971 => (x"00",x"44",x"44",x"44"),
  1972 => (x"7c",x"38",x"00",x"00"),
  1973 => (x"7f",x"7f",x"44",x"44"),
  1974 => (x"7c",x"38",x"00",x"00"),
  1975 => (x"18",x"5c",x"54",x"54"),
  1976 => (x"7e",x"04",x"00",x"00"),
  1977 => (x"00",x"05",x"05",x"7f"),
  1978 => (x"bc",x"18",x"00",x"00"),
  1979 => (x"7c",x"fc",x"a4",x"a4"),
  1980 => (x"7f",x"7f",x"00",x"00"),
  1981 => (x"78",x"7c",x"04",x"04"),
  1982 => (x"00",x"00",x"00",x"00"),
  1983 => (x"00",x"40",x"7d",x"3d"),
  1984 => (x"80",x"80",x"00",x"00"),
  1985 => (x"00",x"7d",x"fd",x"80"),
  1986 => (x"7f",x"7f",x"00",x"00"),
  1987 => (x"44",x"6c",x"38",x"10"),
  1988 => (x"00",x"00",x"00",x"00"),
  1989 => (x"00",x"40",x"7f",x"3f"),
  1990 => (x"0c",x"7c",x"7c",x"00"),
  1991 => (x"78",x"7c",x"0c",x"18"),
  1992 => (x"7c",x"7c",x"00",x"00"),
  1993 => (x"78",x"7c",x"04",x"04"),
  1994 => (x"7c",x"38",x"00",x"00"),
  1995 => (x"38",x"7c",x"44",x"44"),
  1996 => (x"fc",x"fc",x"00",x"00"),
  1997 => (x"18",x"3c",x"24",x"24"),
  1998 => (x"3c",x"18",x"00",x"00"),
  1999 => (x"fc",x"fc",x"24",x"24"),
  2000 => (x"7c",x"7c",x"00",x"00"),
  2001 => (x"08",x"0c",x"04",x"04"),
  2002 => (x"5c",x"48",x"00",x"00"),
  2003 => (x"20",x"74",x"54",x"54"),
  2004 => (x"3f",x"04",x"00",x"00"),
  2005 => (x"00",x"44",x"44",x"7f"),
  2006 => (x"7c",x"3c",x"00",x"00"),
  2007 => (x"7c",x"7c",x"40",x"40"),
  2008 => (x"3c",x"1c",x"00",x"00"),
  2009 => (x"1c",x"3c",x"60",x"60"),
  2010 => (x"60",x"7c",x"3c",x"00"),
  2011 => (x"3c",x"7c",x"60",x"30"),
  2012 => (x"38",x"6c",x"44",x"00"),
  2013 => (x"44",x"6c",x"38",x"10"),
  2014 => (x"bc",x"1c",x"00",x"00"),
  2015 => (x"1c",x"3c",x"60",x"e0"),
  2016 => (x"64",x"44",x"00",x"00"),
  2017 => (x"44",x"4c",x"5c",x"74"),
  2018 => (x"08",x"08",x"00",x"00"),
  2019 => (x"41",x"41",x"77",x"3e"),
  2020 => (x"00",x"00",x"00",x"00"),
  2021 => (x"00",x"00",x"7f",x"7f"),
  2022 => (x"41",x"41",x"00",x"00"),
  2023 => (x"08",x"08",x"3e",x"77"),
  2024 => (x"01",x"01",x"02",x"00"),
  2025 => (x"01",x"02",x"02",x"03"),
  2026 => (x"7f",x"7f",x"7f",x"00"),
  2027 => (x"7f",x"7f",x"7f",x"7f"),
  2028 => (x"1c",x"08",x"08",x"00"),
  2029 => (x"7f",x"3e",x"3e",x"1c"),
  2030 => (x"3e",x"7f",x"7f",x"7f"),
  2031 => (x"08",x"1c",x"1c",x"3e"),
  2032 => (x"18",x"10",x"00",x"08"),
  2033 => (x"10",x"18",x"7c",x"7c"),
  2034 => (x"30",x"10",x"00",x"00"),
  2035 => (x"10",x"30",x"7c",x"7c"),
  2036 => (x"60",x"30",x"10",x"00"),
  2037 => (x"06",x"1e",x"78",x"60"),
  2038 => (x"3c",x"66",x"42",x"00"),
  2039 => (x"42",x"66",x"3c",x"18"),
  2040 => (x"6a",x"38",x"78",x"00"),
  2041 => (x"38",x"6c",x"c6",x"c2"),
  2042 => (x"00",x"00",x"60",x"00"),
  2043 => (x"60",x"00",x"00",x"60"),
  2044 => (x"5b",x"5e",x"0e",x"00"),
  2045 => (x"1e",x"0e",x"5d",x"5c"),
  2046 => (x"f4",x"c2",x"4c",x"71"),
  2047 => (x"c0",x"4d",x"bf",x"c9"),
  2048 => (x"74",x"1e",x"c0",x"4b"),
  2049 => (x"87",x"c7",x"02",x"ab"),
  2050 => (x"c0",x"48",x"a6",x"c4"),
  2051 => (x"c4",x"87",x"c5",x"78"),
  2052 => (x"78",x"c1",x"48",x"a6"),
  2053 => (x"73",x"1e",x"66",x"c4"),
  2054 => (x"87",x"df",x"ee",x"49"),
  2055 => (x"e0",x"c0",x"86",x"c8"),
  2056 => (x"87",x"ef",x"ef",x"49"),
  2057 => (x"6a",x"4a",x"a5",x"c4"),
  2058 => (x"87",x"f0",x"f0",x"49"),
  2059 => (x"cb",x"87",x"c6",x"f1"),
  2060 => (x"c8",x"83",x"c1",x"85"),
  2061 => (x"ff",x"04",x"ab",x"b7"),
  2062 => (x"26",x"26",x"87",x"c7"),
  2063 => (x"26",x"4c",x"26",x"4d"),
  2064 => (x"1e",x"4f",x"26",x"4b"),
  2065 => (x"f4",x"c2",x"4a",x"71"),
  2066 => (x"f4",x"c2",x"5a",x"cd"),
  2067 => (x"78",x"c7",x"48",x"cd"),
  2068 => (x"87",x"dd",x"fe",x"49"),
  2069 => (x"73",x"1e",x"4f",x"26"),
  2070 => (x"c0",x"4a",x"71",x"1e"),
  2071 => (x"d3",x"03",x"aa",x"b7"),
  2072 => (x"d3",x"cf",x"c2",x"87"),
  2073 => (x"87",x"c4",x"05",x"bf"),
  2074 => (x"87",x"c2",x"4b",x"c1"),
  2075 => (x"cf",x"c2",x"4b",x"c0"),
  2076 => (x"87",x"c4",x"5b",x"d7"),
  2077 => (x"5a",x"d7",x"cf",x"c2"),
  2078 => (x"bf",x"d3",x"cf",x"c2"),
  2079 => (x"c1",x"9a",x"c1",x"4a"),
  2080 => (x"ec",x"49",x"a2",x"c0"),
  2081 => (x"48",x"fc",x"87",x"e8"),
  2082 => (x"bf",x"d3",x"cf",x"c2"),
  2083 => (x"87",x"ef",x"fe",x"78"),
  2084 => (x"c4",x"4a",x"71",x"1e"),
  2085 => (x"49",x"72",x"1e",x"66"),
  2086 => (x"26",x"87",x"f9",x"ea"),
  2087 => (x"71",x"1e",x"4f",x"26"),
  2088 => (x"48",x"d4",x"ff",x"4a"),
  2089 => (x"ff",x"78",x"ff",x"c3"),
  2090 => (x"e1",x"c0",x"48",x"d0"),
  2091 => (x"48",x"d4",x"ff",x"78"),
  2092 => (x"49",x"72",x"78",x"c1"),
  2093 => (x"78",x"71",x"31",x"c4"),
  2094 => (x"c0",x"48",x"d0",x"ff"),
  2095 => (x"4f",x"26",x"78",x"e0"),
  2096 => (x"d3",x"cf",x"c2",x"1e"),
  2097 => (x"cb",x"da",x"49",x"bf"),
  2098 => (x"c1",x"f4",x"c2",x"87"),
  2099 => (x"78",x"bf",x"e8",x"48"),
  2100 => (x"48",x"fd",x"f3",x"c2"),
  2101 => (x"c2",x"78",x"bf",x"ec"),
  2102 => (x"4a",x"bf",x"c1",x"f4"),
  2103 => (x"99",x"ff",x"c3",x"49"),
  2104 => (x"72",x"2a",x"b7",x"c8"),
  2105 => (x"c2",x"b0",x"71",x"48"),
  2106 => (x"26",x"58",x"c9",x"f4"),
  2107 => (x"5b",x"5e",x"0e",x"4f"),
  2108 => (x"71",x"0e",x"5d",x"5c"),
  2109 => (x"87",x"c8",x"ff",x"4b"),
  2110 => (x"48",x"fc",x"f3",x"c2"),
  2111 => (x"49",x"73",x"50",x"c0"),
  2112 => (x"70",x"87",x"ee",x"e6"),
  2113 => (x"9c",x"c2",x"4c",x"49"),
  2114 => (x"cb",x"49",x"ee",x"cb"),
  2115 => (x"49",x"70",x"87",x"cd"),
  2116 => (x"fc",x"f3",x"c2",x"4d"),
  2117 => (x"c1",x"05",x"bf",x"97"),
  2118 => (x"66",x"d0",x"87",x"e2"),
  2119 => (x"c5",x"f4",x"c2",x"49"),
  2120 => (x"d6",x"05",x"99",x"bf"),
  2121 => (x"49",x"66",x"d4",x"87"),
  2122 => (x"bf",x"fd",x"f3",x"c2"),
  2123 => (x"87",x"cb",x"05",x"99"),
  2124 => (x"fc",x"e5",x"49",x"73"),
  2125 => (x"02",x"98",x"70",x"87"),
  2126 => (x"c1",x"87",x"c1",x"c1"),
  2127 => (x"87",x"c0",x"fe",x"4c"),
  2128 => (x"e2",x"ca",x"49",x"75"),
  2129 => (x"02",x"98",x"70",x"87"),
  2130 => (x"f3",x"c2",x"87",x"c6"),
  2131 => (x"50",x"c1",x"48",x"fc"),
  2132 => (x"97",x"fc",x"f3",x"c2"),
  2133 => (x"e3",x"c0",x"05",x"bf"),
  2134 => (x"c5",x"f4",x"c2",x"87"),
  2135 => (x"66",x"d0",x"49",x"bf"),
  2136 => (x"d6",x"ff",x"05",x"99"),
  2137 => (x"fd",x"f3",x"c2",x"87"),
  2138 => (x"66",x"d4",x"49",x"bf"),
  2139 => (x"ca",x"ff",x"05",x"99"),
  2140 => (x"e4",x"49",x"73",x"87"),
  2141 => (x"98",x"70",x"87",x"fb"),
  2142 => (x"87",x"ff",x"fe",x"05"),
  2143 => (x"fa",x"fa",x"48",x"74"),
  2144 => (x"5b",x"5e",x"0e",x"87"),
  2145 => (x"f8",x"0e",x"5d",x"5c"),
  2146 => (x"4c",x"4d",x"c0",x"86"),
  2147 => (x"c4",x"7e",x"bf",x"ec"),
  2148 => (x"f4",x"c2",x"48",x"a6"),
  2149 => (x"c1",x"78",x"bf",x"c9"),
  2150 => (x"c7",x"1e",x"c0",x"1e"),
  2151 => (x"87",x"cd",x"fd",x"49"),
  2152 => (x"98",x"70",x"86",x"c8"),
  2153 => (x"ff",x"87",x"cd",x"02"),
  2154 => (x"87",x"ea",x"fa",x"49"),
  2155 => (x"e3",x"49",x"da",x"c1"),
  2156 => (x"4d",x"c1",x"87",x"ff"),
  2157 => (x"97",x"fc",x"f3",x"c2"),
  2158 => (x"87",x"cf",x"02",x"bf"),
  2159 => (x"bf",x"cb",x"cf",x"c2"),
  2160 => (x"c2",x"b9",x"c1",x"49"),
  2161 => (x"71",x"59",x"cf",x"cf"),
  2162 => (x"c2",x"87",x"d3",x"fb"),
  2163 => (x"4b",x"bf",x"c1",x"f4"),
  2164 => (x"bf",x"d3",x"cf",x"c2"),
  2165 => (x"87",x"e9",x"c0",x"05"),
  2166 => (x"e3",x"49",x"fd",x"c3"),
  2167 => (x"fa",x"c3",x"87",x"d3"),
  2168 => (x"87",x"cd",x"e3",x"49"),
  2169 => (x"ff",x"c3",x"49",x"73"),
  2170 => (x"c0",x"1e",x"71",x"99"),
  2171 => (x"87",x"e0",x"fa",x"49"),
  2172 => (x"b7",x"c8",x"49",x"73"),
  2173 => (x"c1",x"1e",x"71",x"29"),
  2174 => (x"87",x"d4",x"fa",x"49"),
  2175 => (x"f4",x"c5",x"86",x"c8"),
  2176 => (x"c5",x"f4",x"c2",x"87"),
  2177 => (x"02",x"9b",x"4b",x"bf"),
  2178 => (x"cf",x"c2",x"87",x"dd"),
  2179 => (x"c7",x"49",x"bf",x"cf"),
  2180 => (x"98",x"70",x"87",x"d5"),
  2181 => (x"c0",x"87",x"c4",x"05"),
  2182 => (x"c2",x"87",x"d2",x"4b"),
  2183 => (x"fa",x"c6",x"49",x"e0"),
  2184 => (x"d3",x"cf",x"c2",x"87"),
  2185 => (x"c2",x"87",x"c6",x"58"),
  2186 => (x"c0",x"48",x"cf",x"cf"),
  2187 => (x"c2",x"49",x"73",x"78"),
  2188 => (x"87",x"cd",x"05",x"99"),
  2189 => (x"e1",x"49",x"eb",x"c3"),
  2190 => (x"49",x"70",x"87",x"f7"),
  2191 => (x"c2",x"02",x"99",x"c2"),
  2192 => (x"73",x"4c",x"fb",x"87"),
  2193 => (x"05",x"99",x"c1",x"49"),
  2194 => (x"f4",x"c3",x"87",x"cd"),
  2195 => (x"87",x"e1",x"e1",x"49"),
  2196 => (x"99",x"c2",x"49",x"70"),
  2197 => (x"fa",x"87",x"c2",x"02"),
  2198 => (x"c8",x"49",x"73",x"4c"),
  2199 => (x"87",x"cd",x"05",x"99"),
  2200 => (x"e1",x"49",x"f5",x"c3"),
  2201 => (x"49",x"70",x"87",x"cb"),
  2202 => (x"d5",x"02",x"99",x"c2"),
  2203 => (x"cd",x"f4",x"c2",x"87"),
  2204 => (x"87",x"ca",x"02",x"bf"),
  2205 => (x"c2",x"88",x"c1",x"48"),
  2206 => (x"c0",x"58",x"d1",x"f4"),
  2207 => (x"4c",x"ff",x"87",x"c2"),
  2208 => (x"49",x"73",x"4d",x"c1"),
  2209 => (x"cd",x"05",x"99",x"c4"),
  2210 => (x"49",x"f2",x"c3",x"87"),
  2211 => (x"70",x"87",x"e2",x"e0"),
  2212 => (x"02",x"99",x"c2",x"49"),
  2213 => (x"f4",x"c2",x"87",x"dc"),
  2214 => (x"48",x"7e",x"bf",x"cd"),
  2215 => (x"03",x"a8",x"b7",x"c7"),
  2216 => (x"6e",x"87",x"cb",x"c0"),
  2217 => (x"c2",x"80",x"c1",x"48"),
  2218 => (x"c0",x"58",x"d1",x"f4"),
  2219 => (x"4c",x"fe",x"87",x"c2"),
  2220 => (x"fd",x"c3",x"4d",x"c1"),
  2221 => (x"f8",x"df",x"ff",x"49"),
  2222 => (x"c2",x"49",x"70",x"87"),
  2223 => (x"87",x"d5",x"02",x"99"),
  2224 => (x"bf",x"cd",x"f4",x"c2"),
  2225 => (x"87",x"c9",x"c0",x"02"),
  2226 => (x"48",x"cd",x"f4",x"c2"),
  2227 => (x"c2",x"c0",x"78",x"c0"),
  2228 => (x"c1",x"4c",x"fd",x"87"),
  2229 => (x"49",x"fa",x"c3",x"4d"),
  2230 => (x"87",x"d5",x"df",x"ff"),
  2231 => (x"99",x"c2",x"49",x"70"),
  2232 => (x"87",x"d9",x"c0",x"02"),
  2233 => (x"bf",x"cd",x"f4",x"c2"),
  2234 => (x"a8",x"b7",x"c7",x"48"),
  2235 => (x"87",x"c9",x"c0",x"03"),
  2236 => (x"48",x"cd",x"f4",x"c2"),
  2237 => (x"c2",x"c0",x"78",x"c7"),
  2238 => (x"c1",x"4c",x"fc",x"87"),
  2239 => (x"ac",x"b7",x"c0",x"4d"),
  2240 => (x"87",x"d3",x"c0",x"03"),
  2241 => (x"c1",x"48",x"66",x"c4"),
  2242 => (x"7e",x"70",x"80",x"d8"),
  2243 => (x"c0",x"02",x"bf",x"6e"),
  2244 => (x"74",x"4b",x"87",x"c5"),
  2245 => (x"c0",x"0f",x"73",x"49"),
  2246 => (x"1e",x"f0",x"c3",x"1e"),
  2247 => (x"f7",x"49",x"da",x"c1"),
  2248 => (x"86",x"c8",x"87",x"cb"),
  2249 => (x"c0",x"02",x"98",x"70"),
  2250 => (x"f4",x"c2",x"87",x"d8"),
  2251 => (x"6e",x"7e",x"bf",x"cd"),
  2252 => (x"c4",x"91",x"cb",x"49"),
  2253 => (x"82",x"71",x"4a",x"66"),
  2254 => (x"c5",x"c0",x"02",x"6a"),
  2255 => (x"49",x"6e",x"4b",x"87"),
  2256 => (x"9d",x"75",x"0f",x"73"),
  2257 => (x"87",x"c8",x"c0",x"02"),
  2258 => (x"bf",x"cd",x"f4",x"c2"),
  2259 => (x"87",x"e1",x"f2",x"49"),
  2260 => (x"bf",x"d7",x"cf",x"c2"),
  2261 => (x"87",x"dd",x"c0",x"02"),
  2262 => (x"87",x"cb",x"c2",x"49"),
  2263 => (x"c0",x"02",x"98",x"70"),
  2264 => (x"f4",x"c2",x"87",x"d3"),
  2265 => (x"f2",x"49",x"bf",x"cd"),
  2266 => (x"49",x"c0",x"87",x"c7"),
  2267 => (x"c2",x"87",x"e7",x"f3"),
  2268 => (x"c0",x"48",x"d7",x"cf"),
  2269 => (x"f3",x"8e",x"f8",x"78"),
  2270 => (x"5e",x"0e",x"87",x"c1"),
  2271 => (x"0e",x"5d",x"5c",x"5b"),
  2272 => (x"c2",x"4c",x"71",x"1e"),
  2273 => (x"49",x"bf",x"c9",x"f4"),
  2274 => (x"4d",x"a1",x"cd",x"c1"),
  2275 => (x"69",x"81",x"d1",x"c1"),
  2276 => (x"02",x"9c",x"74",x"7e"),
  2277 => (x"a5",x"c4",x"87",x"cf"),
  2278 => (x"c2",x"7b",x"74",x"4b"),
  2279 => (x"49",x"bf",x"c9",x"f4"),
  2280 => (x"6e",x"87",x"e0",x"f2"),
  2281 => (x"05",x"9c",x"74",x"7b"),
  2282 => (x"4b",x"c0",x"87",x"c4"),
  2283 => (x"4b",x"c1",x"87",x"c2"),
  2284 => (x"e1",x"f2",x"49",x"73"),
  2285 => (x"02",x"66",x"d4",x"87"),
  2286 => (x"de",x"49",x"87",x"c7"),
  2287 => (x"c2",x"4a",x"70",x"87"),
  2288 => (x"c2",x"4a",x"c0",x"87"),
  2289 => (x"26",x"5a",x"db",x"cf"),
  2290 => (x"00",x"87",x"f0",x"f1"),
  2291 => (x"00",x"00",x"00",x"00"),
  2292 => (x"00",x"00",x"00",x"00"),
  2293 => (x"00",x"00",x"00",x"00"),
  2294 => (x"1e",x"00",x"00",x"00"),
  2295 => (x"c8",x"ff",x"4a",x"71"),
  2296 => (x"a1",x"72",x"49",x"bf"),
  2297 => (x"1e",x"4f",x"26",x"48"),
  2298 => (x"89",x"bf",x"c8",x"ff"),
  2299 => (x"c0",x"c0",x"c0",x"fe"),
  2300 => (x"01",x"a9",x"c0",x"c0"),
  2301 => (x"4a",x"c0",x"87",x"c4"),
  2302 => (x"4a",x"c1",x"87",x"c2"),
  2303 => (x"4f",x"26",x"48",x"72"),
  2304 => (x"dc",x"d3",x"ff",x"1e"),
  2305 => (x"49",x"66",x"c4",x"87"),
  2306 => (x"02",x"99",x"c0",x"c2"),
  2307 => (x"e0",x"c3",x"87",x"cd"),
  2308 => (x"de",x"f3",x"c2",x"1e"),
  2309 => (x"eb",x"d4",x"ff",x"49"),
  2310 => (x"c4",x"86",x"c4",x"87"),
  2311 => (x"c0",x"c4",x"49",x"66"),
  2312 => (x"87",x"cd",x"02",x"99"),
  2313 => (x"c2",x"1e",x"f0",x"c3"),
  2314 => (x"ff",x"49",x"de",x"f3"),
  2315 => (x"c4",x"87",x"d5",x"d4"),
  2316 => (x"49",x"66",x"c4",x"86"),
  2317 => (x"71",x"99",x"ff",x"c1"),
  2318 => (x"de",x"f3",x"c2",x"1e"),
  2319 => (x"c3",x"d4",x"ff",x"49"),
  2320 => (x"d4",x"d2",x"ff",x"87"),
  2321 => (x"4f",x"26",x"26",x"87"),
  2322 => (x"5c",x"5b",x"5e",x"0e"),
  2323 => (x"dc",x"ff",x"0e",x"5d"),
  2324 => (x"c2",x"7e",x"c0",x"86"),
  2325 => (x"49",x"bf",x"d5",x"f4"),
  2326 => (x"1e",x"71",x"81",x"c2"),
  2327 => (x"4a",x"c6",x"1e",x"72"),
  2328 => (x"87",x"c7",x"f2",x"fd"),
  2329 => (x"4a",x"26",x"48",x"71"),
  2330 => (x"a6",x"c8",x"49",x"26"),
  2331 => (x"d5",x"f4",x"c2",x"58"),
  2332 => (x"81",x"c4",x"49",x"bf"),
  2333 => (x"1e",x"72",x"1e",x"71"),
  2334 => (x"f1",x"fd",x"4a",x"c6"),
  2335 => (x"48",x"71",x"87",x"ed"),
  2336 => (x"49",x"26",x"4a",x"26"),
  2337 => (x"c2",x"58",x"a6",x"cc"),
  2338 => (x"49",x"bf",x"ee",x"dc"),
  2339 => (x"70",x"87",x"d8",x"fd"),
  2340 => (x"ce",x"ca",x"02",x"98"),
  2341 => (x"49",x"e0",x"c0",x"87"),
  2342 => (x"70",x"87",x"c0",x"fd"),
  2343 => (x"f2",x"dc",x"c2",x"49"),
  2344 => (x"74",x"4c",x"c0",x"59"),
  2345 => (x"fe",x"91",x"c4",x"49"),
  2346 => (x"4a",x"69",x"81",x"d0"),
  2347 => (x"f4",x"c2",x"49",x"74"),
  2348 => (x"c4",x"81",x"bf",x"d5"),
  2349 => (x"e5",x"f4",x"c2",x"91"),
  2350 => (x"9a",x"79",x"72",x"81"),
  2351 => (x"72",x"87",x"d2",x"02"),
  2352 => (x"71",x"89",x"c1",x"49"),
  2353 => (x"c1",x"48",x"6e",x"9a"),
  2354 => (x"72",x"7e",x"70",x"80"),
  2355 => (x"ee",x"ff",x"05",x"9a"),
  2356 => (x"c2",x"84",x"c1",x"87"),
  2357 => (x"ff",x"04",x"ac",x"b7"),
  2358 => (x"48",x"6e",x"87",x"c9"),
  2359 => (x"a8",x"b7",x"fc",x"c0"),
  2360 => (x"87",x"ff",x"c8",x"04"),
  2361 => (x"4a",x"74",x"4c",x"c0"),
  2362 => (x"c4",x"82",x"66",x"c4"),
  2363 => (x"e5",x"f4",x"c2",x"92"),
  2364 => (x"c8",x"49",x"74",x"82"),
  2365 => (x"91",x"c4",x"81",x"66"),
  2366 => (x"81",x"e5",x"f4",x"c2"),
  2367 => (x"49",x"69",x"4a",x"6a"),
  2368 => (x"4b",x"74",x"b9",x"72"),
  2369 => (x"bf",x"d5",x"f4",x"c2"),
  2370 => (x"c2",x"93",x"c4",x"83"),
  2371 => (x"6b",x"83",x"e5",x"f4"),
  2372 => (x"71",x"48",x"72",x"ba"),
  2373 => (x"58",x"a6",x"d0",x"98"),
  2374 => (x"f4",x"c2",x"49",x"74"),
  2375 => (x"c4",x"81",x"bf",x"d5"),
  2376 => (x"e5",x"f4",x"c2",x"91"),
  2377 => (x"d0",x"7e",x"69",x"81"),
  2378 => (x"78",x"c0",x"48",x"a6"),
  2379 => (x"df",x"49",x"66",x"cc"),
  2380 => (x"c0",x"c7",x"02",x"29"),
  2381 => (x"c0",x"4a",x"74",x"87"),
  2382 => (x"66",x"d0",x"92",x"e0"),
  2383 => (x"48",x"ff",x"c0",x"82"),
  2384 => (x"4a",x"70",x"88",x"72"),
  2385 => (x"c0",x"48",x"a6",x"d4"),
  2386 => (x"c0",x"80",x"c4",x"78"),
  2387 => (x"df",x"49",x"6e",x"78"),
  2388 => (x"a6",x"e0",x"c0",x"29"),
  2389 => (x"d1",x"f4",x"c2",x"59"),
  2390 => (x"72",x"78",x"c1",x"48"),
  2391 => (x"b7",x"31",x"c3",x"49"),
  2392 => (x"c0",x"b1",x"72",x"2a"),
  2393 => (x"91",x"c4",x"99",x"ff"),
  2394 => (x"4d",x"c5",x"de",x"c2"),
  2395 => (x"4b",x"6d",x"85",x"71"),
  2396 => (x"c0",x"c0",x"c4",x"49"),
  2397 => (x"f3",x"c0",x"02",x"99"),
  2398 => (x"02",x"66",x"dc",x"87"),
  2399 => (x"80",x"c8",x"87",x"c8"),
  2400 => (x"c5",x"78",x"40",x"c0"),
  2401 => (x"f4",x"c2",x"87",x"ef"),
  2402 => (x"78",x"c1",x"48",x"d9"),
  2403 => (x"bf",x"dd",x"f4",x"c2"),
  2404 => (x"87",x"e1",x"c5",x"05"),
  2405 => (x"f8",x"1e",x"d8",x"c1"),
  2406 => (x"e3",x"f9",x"49",x"a0"),
  2407 => (x"1e",x"d8",x"c5",x"87"),
  2408 => (x"49",x"d1",x"f4",x"c2"),
  2409 => (x"c8",x"87",x"d9",x"f9"),
  2410 => (x"87",x"c9",x"c5",x"86"),
  2411 => (x"d8",x"02",x"66",x"dc"),
  2412 => (x"c2",x"49",x"73",x"87"),
  2413 => (x"02",x"99",x"c0",x"c0"),
  2414 => (x"d0",x"87",x"c3",x"c0"),
  2415 => (x"48",x"6d",x"2b",x"b7"),
  2416 => (x"98",x"ff",x"ff",x"fd"),
  2417 => (x"fa",x"c0",x"7d",x"70"),
  2418 => (x"d9",x"f4",x"c2",x"87"),
  2419 => (x"f2",x"c0",x"02",x"bf"),
  2420 => (x"d0",x"48",x"73",x"87"),
  2421 => (x"e4",x"c0",x"28",x"b7"),
  2422 => (x"98",x"70",x"58",x"a6"),
  2423 => (x"87",x"e3",x"c0",x"02"),
  2424 => (x"bf",x"e1",x"f4",x"c2"),
  2425 => (x"c0",x"e0",x"c0",x"49"),
  2426 => (x"ca",x"c0",x"02",x"99"),
  2427 => (x"c0",x"49",x"70",x"87"),
  2428 => (x"02",x"99",x"c0",x"e0"),
  2429 => (x"6d",x"87",x"cc",x"c0"),
  2430 => (x"c0",x"c0",x"c2",x"48"),
  2431 => (x"c0",x"7d",x"70",x"b0"),
  2432 => (x"73",x"4b",x"66",x"e0"),
  2433 => (x"c0",x"c0",x"c8",x"49"),
  2434 => (x"c7",x"c2",x"02",x"99"),
  2435 => (x"e1",x"f4",x"c2",x"87"),
  2436 => (x"c0",x"cc",x"4a",x"bf"),
  2437 => (x"cf",x"c0",x"02",x"9a"),
  2438 => (x"8a",x"c0",x"c4",x"87"),
  2439 => (x"87",x"d8",x"c0",x"02"),
  2440 => (x"f9",x"c0",x"02",x"8a"),
  2441 => (x"87",x"dd",x"c1",x"87"),
  2442 => (x"ff",x"c3",x"49",x"73"),
  2443 => (x"c2",x"91",x"c2",x"99"),
  2444 => (x"11",x"81",x"f9",x"dd"),
  2445 => (x"87",x"dc",x"c1",x"4b"),
  2446 => (x"ff",x"c3",x"49",x"73"),
  2447 => (x"c2",x"91",x"c2",x"99"),
  2448 => (x"c1",x"81",x"f9",x"dd"),
  2449 => (x"dc",x"4b",x"11",x"81"),
  2450 => (x"c8",x"c0",x"02",x"66"),
  2451 => (x"48",x"a6",x"d8",x"87"),
  2452 => (x"ff",x"c0",x"78",x"d2"),
  2453 => (x"48",x"a6",x"d4",x"87"),
  2454 => (x"c0",x"78",x"d2",x"c4"),
  2455 => (x"49",x"73",x"87",x"f6"),
  2456 => (x"c2",x"99",x"ff",x"c3"),
  2457 => (x"f9",x"dd",x"c2",x"91"),
  2458 => (x"11",x"81",x"c1",x"81"),
  2459 => (x"02",x"66",x"dc",x"4b"),
  2460 => (x"d8",x"87",x"c9",x"c0"),
  2461 => (x"d9",x"c1",x"48",x"a6"),
  2462 => (x"87",x"d8",x"c0",x"78"),
  2463 => (x"c5",x"48",x"a6",x"d4"),
  2464 => (x"cf",x"c0",x"78",x"d9"),
  2465 => (x"c3",x"49",x"73",x"87"),
  2466 => (x"91",x"c2",x"99",x"ff"),
  2467 => (x"81",x"f9",x"dd",x"c2"),
  2468 => (x"4b",x"11",x"81",x"c1"),
  2469 => (x"c0",x"02",x"66",x"dc"),
  2470 => (x"49",x"73",x"87",x"dc"),
  2471 => (x"fc",x"c7",x"b9",x"ff"),
  2472 => (x"48",x"71",x"99",x"c0"),
  2473 => (x"bf",x"e1",x"f4",x"c2"),
  2474 => (x"e5",x"f4",x"c2",x"98"),
  2475 => (x"9b",x"ff",x"c3",x"58"),
  2476 => (x"c0",x"b3",x"c0",x"c4"),
  2477 => (x"49",x"73",x"87",x"d4"),
  2478 => (x"99",x"c0",x"fc",x"c7"),
  2479 => (x"f4",x"c2",x"48",x"71"),
  2480 => (x"c2",x"b0",x"bf",x"e1"),
  2481 => (x"c3",x"58",x"e5",x"f4"),
  2482 => (x"66",x"d4",x"9b",x"ff"),
  2483 => (x"87",x"ca",x"c0",x"02"),
  2484 => (x"d1",x"f4",x"c2",x"1e"),
  2485 => (x"87",x"e8",x"f4",x"49"),
  2486 => (x"1e",x"73",x"86",x"c4"),
  2487 => (x"49",x"d1",x"f4",x"c2"),
  2488 => (x"c4",x"87",x"dd",x"f4"),
  2489 => (x"02",x"66",x"d8",x"86"),
  2490 => (x"1e",x"87",x"ca",x"c0"),
  2491 => (x"49",x"d1",x"f4",x"c2"),
  2492 => (x"c4",x"87",x"cd",x"f4"),
  2493 => (x"48",x"66",x"cc",x"86"),
  2494 => (x"a6",x"d0",x"30",x"c1"),
  2495 => (x"c1",x"48",x"6e",x"58"),
  2496 => (x"d0",x"7e",x"70",x"30"),
  2497 => (x"80",x"c1",x"48",x"66"),
  2498 => (x"c0",x"58",x"a6",x"d4"),
  2499 => (x"04",x"a8",x"b7",x"e0"),
  2500 => (x"c1",x"87",x"d9",x"f8"),
  2501 => (x"ac",x"b7",x"c2",x"84"),
  2502 => (x"87",x"ca",x"f7",x"04"),
  2503 => (x"48",x"d5",x"f4",x"c2"),
  2504 => (x"ff",x"78",x"66",x"c4"),
  2505 => (x"4d",x"26",x"8e",x"dc"),
  2506 => (x"4b",x"26",x"4c",x"26"),
  2507 => (x"00",x"00",x"4f",x"26"),
  2508 => (x"c0",x"1e",x"00",x"00"),
  2509 => (x"c4",x"49",x"72",x"4a"),
  2510 => (x"e5",x"f4",x"c2",x"91"),
  2511 => (x"c1",x"79",x"ff",x"81"),
  2512 => (x"aa",x"b7",x"c6",x"82"),
  2513 => (x"c2",x"87",x"ee",x"04"),
  2514 => (x"c0",x"48",x"d5",x"f4"),
  2515 => (x"80",x"c8",x"78",x"40"),
  2516 => (x"4f",x"26",x"78",x"c0"),
  2517 => (x"71",x"1e",x"73",x"1e"),
  2518 => (x"f5",x"dd",x"c2",x"4b"),
  2519 => (x"87",x"c9",x"05",x"bf"),
  2520 => (x"48",x"f5",x"dd",x"c2"),
  2521 => (x"c9",x"ff",x"78",x"c1"),
  2522 => (x"87",x"dc",x"f3",x"87"),
  2523 => (x"c8",x"ff",x"49",x"73"),
  2524 => (x"f5",x"fe",x"87",x"fc"),
  2525 => (x"00",x"00",x"00",x"87"),
  2526 => (x"f2",x"eb",x"f4",x"00"),
  2527 => (x"04",x"06",x"05",x"f5"),
  2528 => (x"83",x"0b",x"03",x"0c"),
  2529 => (x"fc",x"00",x"66",x"0a"),
  2530 => (x"da",x"00",x"5a",x"00"),
  2531 => (x"94",x"80",x"00",x"00"),
  2532 => (x"78",x"80",x"05",x"08"),
  2533 => (x"01",x"80",x"02",x"00"),
  2534 => (x"09",x"80",x"03",x"00"),
  2535 => (x"00",x"80",x"04",x"00"),
  2536 => (x"91",x"80",x"01",x"00"),
  2537 => (x"04",x"00",x"26",x"08"),
  2538 => (x"00",x"00",x"1d",x"00"),
  2539 => (x"00",x"00",x"1c",x"00"),
  2540 => (x"0c",x"00",x"25",x"00"),
  2541 => (x"00",x"00",x"1a",x"00"),
  2542 => (x"00",x"00",x"1b",x"00"),
  2543 => (x"00",x"00",x"24",x"00"),
  2544 => (x"00",x"01",x"12",x"00"),
  2545 => (x"03",x"00",x"2e",x"00"),
  2546 => (x"00",x"00",x"2d",x"00"),
  2547 => (x"00",x"00",x"23",x"00"),
  2548 => (x"0b",x"00",x"36",x"00"),
  2549 => (x"00",x"00",x"21",x"00"),
  2550 => (x"00",x"00",x"2b",x"00"),
  2551 => (x"00",x"00",x"2c",x"00"),
  2552 => (x"00",x"00",x"22",x"00"),
  2553 => (x"6c",x"00",x"3d",x"00"),
  2554 => (x"00",x"00",x"35",x"00"),
  2555 => (x"00",x"00",x"34",x"00"),
  2556 => (x"75",x"00",x"3e",x"00"),
  2557 => (x"00",x"00",x"32",x"00"),
  2558 => (x"00",x"00",x"33",x"00"),
  2559 => (x"6b",x"00",x"3c",x"00"),
  2560 => (x"00",x"00",x"2a",x"00"),
  2561 => (x"01",x"00",x"46",x"00"),
  2562 => (x"73",x"00",x"43",x"00"),
  2563 => (x"69",x"00",x"3b",x"00"),
  2564 => (x"09",x"00",x"45",x"00"),
  2565 => (x"70",x"00",x"3a",x"00"),
  2566 => (x"72",x"00",x"42",x"00"),
  2567 => (x"74",x"00",x"44",x"00"),
  2568 => (x"00",x"00",x"31",x"00"),
  2569 => (x"00",x"00",x"55",x"00"),
  2570 => (x"7c",x"00",x"4d",x"00"),
  2571 => (x"7a",x"00",x"4b",x"00"),
  2572 => (x"00",x"00",x"7b",x"00"),
  2573 => (x"71",x"00",x"49",x"00"),
  2574 => (x"84",x"00",x"4c",x"00"),
  2575 => (x"77",x"00",x"54",x"00"),
  2576 => (x"00",x"00",x"41",x"00"),
  2577 => (x"00",x"00",x"61",x"00"),
  2578 => (x"7c",x"00",x"5b",x"00"),
  2579 => (x"00",x"00",x"52",x"00"),
  2580 => (x"00",x"00",x"f1",x"00"),
  2581 => (x"00",x"02",x"59",x"00"),
  2582 => (x"5d",x"00",x"0e",x"00"),
  2583 => (x"00",x"00",x"5d",x"00"),
  2584 => (x"79",x"00",x"4a",x"00"),
  2585 => (x"05",x"00",x"16",x"00"),
  2586 => (x"07",x"00",x"76",x"00"),
  2587 => (x"0d",x"00",x"0d",x"00"),
  2588 => (x"06",x"00",x"1e",x"00"),
  2589 => (x"00",x"00",x"29",x"00"),
  2590 => (x"00",x"04",x"14",x"00"),
  2591 => (x"00",x"00",x"15",x"00"),
  2592 => (x"00",x"40",x"00",x"00"),
  2593 => (x"00",x"40",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

